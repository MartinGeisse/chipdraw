magic
tech concept
timestamp 1576406192396
<< sizer >>
rect 0 0 35 140
<< metal1 >>
rect 0 134 35 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 35 134
rect 0 128 35 132
rect 11 124 15 128
rect 19 124 23 125
rect 11 122 12 124
rect 14 122 15 124
rect 19 122 20 124
rect 22 122 23 124
rect 11 120 15 122
rect 19 120 23 122
rect 11 118 12 120
rect 14 118 15 120
rect 19 118 20 120
rect 22 118 23 120
rect 11 117 15 118
rect 19 76 23 118
rect 8 75 17 76
rect 19 72 26 76
rect 8 73 14 75
rect 16 73 17 75
rect 8 72 17 73
rect 19 19 23 72
rect 11 19 15 20
rect 11 17 12 19
rect 14 17 15 19
rect 19 17 20 19
rect 22 17 23 19
rect 11 13 15 17
rect 19 16 23 17
rect 0 8 35 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 35 8
rect 0 2 35 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 12 122 14 124
rect 20 122 22 124
rect 12 118 14 120
rect 20 118 22 120
rect 14 73 16 75
rect 12 17 14 19
rect 20 17 22 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
<< poly >>
rect 16 77 18 128
rect 12 71 18 77
rect 16 13 18 71
<< ndiff >>
rect 6 130 29 136
rect 10 15 24 21
<< pdiff >>
rect 10 116 24 126
rect 6 4 29 10
<< nwell >>
rect 3 48 32 139
<< pwell >>
rect 3 1 32 46
<< end >>
