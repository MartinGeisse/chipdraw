magic
tech concept
timestamp 1577805715535
<< sizer >>
rect 0 0 63 70
<< metal1 >>
rect 0 65 63 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 45 65
rect 47 63 49 65
rect 51 63 53 65
rect 55 63 63 65
rect 0 58 63 63
rect 6 55 14 58
rect 28 50 32 58
rect 36 53 56 56
rect 6 53 7 55
rect 9 53 11 55
rect 13 53 14 55
rect 6 52 14 53
rect 36 50 40 53
rect 52 50 56 53
rect 20 50 24 51
rect 44 50 48 51
rect 20 48 21 50
rect 23 48 24 50
rect 28 48 29 50
rect 31 48 32 50
rect 36 48 37 50
rect 39 48 40 50
rect 44 48 45 50
rect 47 48 48 50
rect 52 48 53 50
rect 55 48 56 50
rect 6 47 14 48
rect 20 46 24 48
rect 28 46 32 48
rect 36 46 40 48
rect 44 46 48 48
rect 52 46 56 48
rect 6 45 7 47
rect 9 45 11 47
rect 13 45 14 47
rect 20 44 21 46
rect 23 44 24 46
rect 28 44 29 46
rect 31 44 32 46
rect 36 44 37 46
rect 39 44 40 46
rect 44 44 45 46
rect 47 44 48 46
rect 52 44 53 46
rect 55 44 56 46
rect 6 44 14 45
rect 11 28 14 44
rect 20 41 24 44
rect 28 43 32 44
rect 36 41 40 44
rect 44 43 48 44
rect 52 43 56 44
rect 45 41 48 43
rect 20 38 40 41
rect 45 38 60 41
rect 57 34 60 38
rect 22 33 26 34
rect 29 33 34 34
rect 42 33 46 34
rect 50 33 54 34
rect 57 30 61 34
rect 22 31 23 33
rect 25 31 26 33
rect 29 31 31 33
rect 33 31 34 33
rect 42 31 43 33
rect 45 31 46 33
rect 50 31 51 33
rect 53 31 54 33
rect 22 30 26 31
rect 29 30 34 31
rect 42 30 46 31
rect 50 30 54 31
rect 42 24 45 30
rect 57 24 60 30
rect 11 25 18 28
rect 15 24 18 25
rect 15 21 45 24
rect 47 21 60 24
rect 15 19 18 21
rect 47 19 50 21
rect 6 18 10 19
rect 14 18 18 19
rect 28 18 32 19
rect 40 18 50 19
rect 52 18 56 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 28 16 29 18
rect 31 16 32 18
rect 40 16 41 18
rect 43 16 50 18
rect 52 16 53 18
rect 55 16 56 18
rect 6 13 10 16
rect 14 15 18 16
rect 28 13 32 16
rect 40 15 44 16
rect 52 13 56 16
rect 0 7 63 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 45 7
rect 47 5 49 7
rect 51 5 53 7
rect 55 5 63 7
rect 0 2 63 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 45 63 47 65
rect 49 63 51 65
rect 53 63 55 65
rect 7 53 9 55
rect 11 53 13 55
rect 21 48 23 50
rect 29 48 31 50
rect 37 48 39 50
rect 45 48 47 50
rect 53 48 55 50
rect 7 45 9 47
rect 11 45 13 47
rect 21 44 23 46
rect 29 44 31 46
rect 37 44 39 46
rect 45 44 47 46
rect 53 44 55 46
rect 23 31 25 33
rect 31 31 33 33
rect 43 31 45 33
rect 51 31 53 33
rect 7 16 9 18
rect 15 16 17 18
rect 29 16 31 18
rect 41 16 43 18
rect 53 16 55 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
rect 45 5 47 7
rect 49 5 51 7
rect 53 5 55 7
<< poly >>
rect 25 41 27 54
rect 33 35 35 54
rect 41 35 43 54
rect 49 35 51 54
rect 3 49 18 51
rect 16 41 18 49
rect 16 39 27 41
rect 21 35 23 39
rect 21 29 27 35
rect 29 31 35 35
rect 41 29 47 35
rect 49 29 56 35
rect 29 29 39 31
rect 21 27 23 29
rect 37 12 39 29
rect 45 12 47 29
rect 49 12 51 29
rect 11 25 35 27
rect 11 12 13 25
rect 33 12 35 25
<< ndiff >>
rect 3 61 60 67
rect 5 14 19 20
rect 27 14 57 20
<< pdiff >>
rect 5 43 15 57
rect 19 42 57 52
rect 3 3 60 9
<< nwell >>
rect 0 31 63 70
<< pwell >>
rect 0 0 63 31
<< end >>
