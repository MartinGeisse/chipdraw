magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577893372126
<< sizer >>
rect 0 0 56 70
<< metal2 >>
rect 26 51 30 52
rect 26 49 27 51
rect 29 49 30 51
rect 26 18 30 49
rect 26 16 27 18
rect 29 16 30 18
rect 26 15 30 16
<< via12 >>
rect 27 49 29 51
rect 27 16 29 18
<< metal1 >>
rect 0 65 56 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 45 65
rect 47 63 49 65
rect 51 63 56 65
rect 0 58 56 63
rect 14 55 18 58
rect 38 55 42 58
rect 6 55 10 56
rect 26 55 30 56
rect 46 55 50 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 26 53 27 55
rect 29 53 30 55
rect 38 53 39 55
rect 41 53 42 55
rect 46 53 47 55
rect 49 53 50 55
rect 6 51 10 53
rect 14 51 18 53
rect 26 51 30 53
rect 38 51 42 53
rect 46 51 50 53
rect 1 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 26 49 27 51
rect 29 49 34 51
rect 38 49 39 51
rect 41 49 42 51
rect 46 49 47 51
rect 49 49 50 51
rect 1 48 10 49
rect 14 48 18 49
rect 26 48 34 49
rect 38 48 42 49
rect 46 48 50 49
rect 1 19 4 48
rect 31 39 34 48
rect 46 46 49 48
rect 8 44 28 46
rect 36 44 53 46
rect 8 42 9 44
rect 11 43 25 44
rect 27 42 28 44
rect 36 42 37 44
rect 39 43 53 44
rect 11 42 12 43
rect 24 42 25 43
rect 39 42 40 43
rect 50 34 53 43
rect 8 41 12 42
rect 24 41 28 42
rect 36 41 40 42
rect 44 40 48 41
rect 44 39 45 40
rect 47 38 48 40
rect 31 38 45 39
rect 31 36 48 38
rect 15 33 19 34
rect 50 30 54 34
rect 15 31 16 33
rect 18 31 19 33
rect 15 30 19 31
rect 50 24 53 30
rect 29 26 32 27
rect 8 25 12 26
rect 28 25 32 26
rect 36 25 40 26
rect 8 23 9 25
rect 11 24 12 25
rect 28 24 29 25
rect 31 23 32 25
rect 36 23 37 25
rect 39 24 40 25
rect 11 23 29 24
rect 39 23 53 24
rect 8 21 32 23
rect 36 21 53 23
rect 46 19 49 21
rect 1 18 10 19
rect 14 18 18 19
rect 26 18 30 19
rect 38 18 42 19
rect 46 18 50 19
rect 1 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 26 16 27 18
rect 29 16 30 18
rect 38 16 39 18
rect 41 16 42 18
rect 46 16 47 18
rect 49 16 50 18
rect 6 15 10 16
rect 14 13 18 16
rect 26 15 30 16
rect 38 13 42 16
rect 46 15 50 16
rect 0 7 56 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 45 7
rect 47 5 49 7
rect 51 5 56 7
rect 0 2 56 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 45 63 47 65
rect 49 63 51 65
rect 7 53 9 55
rect 15 53 17 55
rect 27 53 29 55
rect 39 53 41 55
rect 47 53 49 55
rect 7 49 9 51
rect 15 49 17 51
rect 27 49 29 51
rect 39 49 41 51
rect 47 49 49 51
rect 9 42 11 44
rect 25 42 27 44
rect 37 42 39 44
rect 45 38 47 40
rect 16 31 18 33
rect 9 23 11 25
rect 29 23 31 25
rect 37 23 39 25
rect 7 16 9 18
rect 15 16 17 18
rect 27 16 29 18
rect 39 16 41 18
rect 47 16 49 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
rect 45 5 47 7
rect 49 5 51 7
<< poly >>
rect 11 46 13 59
rect 19 35 21 59
rect 23 46 25 59
rect 31 31 33 59
rect 35 46 37 59
rect 43 42 45 59
rect 7 40 13 46
rect 23 40 29 46
rect 35 40 41 46
rect 43 36 49 42
rect 7 27 9 40
rect 43 12 45 36
rect 14 29 21 35
rect 23 29 33 31
rect 19 12 21 29
rect 23 12 25 29
rect 7 21 13 27
rect 27 21 33 27
rect 35 21 41 27
rect 11 12 13 21
rect 31 12 33 21
rect 35 12 37 21
<< ndiff >>
rect 3 61 53 67
rect 5 14 51 20
<< pdiff >>
rect 5 47 51 57
rect 3 3 53 9
<< nwell >>
rect 0 31 56 70
<< pwell >>
rect 0 0 56 31
<< end >>
