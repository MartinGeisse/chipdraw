magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577092989295
<< sizer >>
rect 0 0 28 70
<< metal1 >>
rect 0 65 28 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 28 65
rect 0 58 28 63
rect 6 55 10 58
rect 18 55 25 56
rect 6 53 7 55
rect 9 53 10 55
rect 18 53 19 55
rect 21 53 25 55
rect 6 51 10 53
rect 18 51 25 53
rect 6 49 7 51
rect 9 49 10 51
rect 18 49 19 51
rect 21 49 25 51
rect 6 48 10 49
rect 18 48 25 49
rect 22 34 25 48
rect 15 40 19 41
rect 15 38 16 40
rect 18 38 19 40
rect 15 37 19 38
rect 1 33 6 34
rect 22 30 26 34
rect 1 31 3 33
rect 5 31 6 33
rect 1 30 6 31
rect 22 19 25 30
rect 15 25 20 27
rect 15 23 17 25
rect 19 23 20 25
rect 15 22 20 23
rect 6 18 10 19
rect 18 18 25 19
rect 6 16 7 18
rect 9 16 10 18
rect 18 16 19 18
rect 21 16 25 18
rect 6 13 10 16
rect 18 15 25 16
rect 0 7 28 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 28 7
rect 0 2 28 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 7 53 9 55
rect 19 53 21 55
rect 7 49 9 51
rect 19 49 21 51
rect 16 38 18 40
rect 3 31 5 33
rect 17 23 19 25
rect 7 16 9 18
rect 19 16 21 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
<< poly >>
rect 11 46 13 59
rect 15 42 17 59
rect 5 44 13 46
rect 5 35 7 44
rect 14 36 20 42
rect 1 29 7 35
rect 5 23 7 29
rect 15 21 21 27
rect 5 21 13 23
rect 11 12 13 21
rect 15 12 17 21
<< ndiff >>
rect 3 61 25 67
rect 5 14 23 20
<< pdiff >>
rect 5 47 23 57
rect 3 3 25 9
<< nwell >>
rect 0 31 28 70
<< pwell >>
rect 0 0 28 31
<< end >>
