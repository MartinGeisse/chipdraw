magic
tech concept
timestamp 1576424724936
<< sizer >>
rect 0 0 42 140
<< metal1 >>
rect 0 134 42 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 28 134
rect 30 132 32 134
rect 34 132 42 134
rect 0 128 42 132
rect 19 124 23 128
rect 10 124 14 125
rect 28 124 32 125
rect 10 122 11 124
rect 13 122 14 124
rect 19 122 20 124
rect 22 122 23 124
rect 28 122 29 124
rect 31 122 32 124
rect 10 120 14 122
rect 19 120 23 122
rect 28 120 32 122
rect 10 118 11 120
rect 13 118 14 120
rect 19 118 20 120
rect 22 118 23 120
rect 28 118 29 120
rect 31 118 32 120
rect 10 117 14 118
rect 19 116 23 118
rect 28 116 32 118
rect 11 90 14 117
rect 19 114 20 116
rect 22 114 23 116
rect 28 114 29 116
rect 31 114 32 116
rect 19 112 23 114
rect 28 112 32 114
rect 19 110 20 112
rect 22 110 23 112
rect 28 110 29 112
rect 31 110 32 112
rect 19 108 23 110
rect 28 76 32 110
rect 19 106 20 108
rect 22 106 23 108
rect 19 104 23 106
rect 19 102 20 104
rect 22 102 23 104
rect 19 100 23 102
rect 19 98 20 100
rect 22 98 23 100
rect 19 96 23 98
rect 19 94 20 96
rect 22 94 23 96
rect 19 93 23 94
rect 11 89 26 90
rect 11 87 23 89
rect 25 87 26 89
rect 22 86 26 87
rect 23 39 26 86
rect 8 75 17 76
rect 28 72 33 76
rect 8 73 14 75
rect 16 73 17 75
rect 8 72 17 73
rect 28 31 32 72
rect 22 38 26 39
rect 11 36 23 38
rect 25 36 26 38
rect 11 35 26 36
rect 11 20 14 35
rect 19 31 23 32
rect 19 29 20 31
rect 22 29 23 31
rect 28 29 29 31
rect 31 29 32 31
rect 19 27 23 29
rect 28 27 32 29
rect 19 25 20 27
rect 22 25 23 27
rect 28 25 29 27
rect 31 25 32 27
rect 19 23 23 25
rect 28 23 32 25
rect 19 21 20 23
rect 22 21 23 23
rect 28 21 29 23
rect 31 21 32 23
rect 19 19 23 21
rect 28 19 32 21
rect 10 19 14 20
rect 10 17 11 19
rect 13 17 14 19
rect 19 17 20 19
rect 22 17 23 19
rect 28 17 29 19
rect 31 17 32 19
rect 10 16 14 17
rect 19 13 23 17
rect 28 16 32 17
rect 0 8 42 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 28 8
rect 30 6 32 8
rect 34 6 42 8
rect 0 2 42 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 28 132 30 134
rect 32 132 34 134
rect 11 122 13 124
rect 20 122 22 124
rect 29 122 31 124
rect 11 118 13 120
rect 20 118 22 120
rect 29 118 31 120
rect 20 114 22 116
rect 29 114 31 116
rect 20 110 22 112
rect 29 110 31 112
rect 20 106 22 108
rect 20 102 22 104
rect 20 98 22 100
rect 20 94 22 96
rect 23 87 25 89
rect 14 73 16 75
rect 23 36 25 38
rect 20 29 22 31
rect 29 29 31 31
rect 20 25 22 27
rect 29 25 31 27
rect 20 21 22 23
rect 29 21 31 23
rect 11 17 13 19
rect 20 17 22 19
rect 29 17 31 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
rect 28 6 30 8
rect 32 6 34 8
<< poly >>
rect 15 77 17 128
rect 25 91 27 128
rect 21 85 27 91
rect 12 71 18 77
rect 15 13 17 71
rect 21 34 27 40
rect 25 13 27 34
<< ndiff >>
rect 6 130 36 136
rect 18 21 33 33
rect 9 15 33 21
<< pdiff >>
rect 9 116 33 126
rect 18 92 33 116
rect 6 4 36 10
<< nwell >>
rect 3 48 39 139
<< pwell >>
rect 3 1 39 46
<< end >>
