magic
tech concept
timestamp 1577800852534
<< sizer >>
rect 0 0 42 70
<< metal1 >>
rect 0 65 42 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 42 65
rect 0 58 42 63
rect 18 55 22 58
rect 6 55 10 56
rect 30 55 34 56
rect 6 53 7 55
rect 9 53 10 55
rect 18 53 19 55
rect 21 53 22 55
rect 30 53 31 55
rect 33 53 34 55
rect 6 51 10 53
rect 18 51 22 53
rect 30 51 34 53
rect 2 49 7 51
rect 9 49 10 51
rect 18 49 19 51
rect 21 49 22 51
rect 30 49 31 51
rect 33 49 39 51
rect 2 48 10 49
rect 18 48 22 49
rect 30 48 39 49
rect 2 34 5 48
rect 36 34 39 48
rect 18 43 22 44
rect 18 41 19 43
rect 21 41 22 43
rect 18 40 22 41
rect 1 30 5 34
rect 7 33 12 34
rect 29 33 33 34
rect 36 30 40 34
rect 7 31 8 33
rect 10 31 12 33
rect 29 31 30 33
rect 32 31 33 33
rect 7 30 12 31
rect 29 30 33 31
rect 2 19 5 30
rect 36 19 39 30
rect 18 26 22 27
rect 18 24 19 26
rect 21 24 22 26
rect 18 23 22 24
rect 2 18 10 19
rect 18 18 22 19
rect 30 18 39 19
rect 2 16 7 18
rect 9 16 10 18
rect 18 16 19 18
rect 21 16 22 18
rect 30 16 31 18
rect 33 16 39 18
rect 6 15 10 16
rect 18 13 22 16
rect 30 15 34 16
rect 0 7 42 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 42 7
rect 0 2 42 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 7 53 9 55
rect 19 53 21 55
rect 31 53 33 55
rect 7 49 9 51
rect 19 49 21 51
rect 31 49 33 51
rect 19 41 21 43
rect 8 31 10 33
rect 30 31 32 33
rect 19 24 21 26
rect 7 16 9 18
rect 19 16 21 18
rect 31 16 33 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
<< poly >>
rect 11 46 13 59
rect 15 45 17 59
rect 23 45 25 59
rect 27 35 29 59
rect 10 44 13 46
rect 15 42 25 45
rect 10 35 12 44
rect 17 39 23 42
rect 6 29 12 35
rect 27 29 34 35
rect 10 23 12 29
rect 27 12 29 29
rect 17 25 23 28
rect 15 22 25 25
rect 10 21 13 23
rect 15 12 17 22
rect 23 12 25 22
rect 11 12 13 21
<< ndiff >>
rect 3 61 39 67
rect 5 14 35 20
<< pdiff >>
rect 5 47 35 57
rect 3 3 39 9
<< nwell >>
rect 0 31 42 70
<< pwell >>
rect 0 0 42 31
<< end >>
