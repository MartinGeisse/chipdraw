magic
tech concept
timestamp 1577173829017
<< sizer >>
rect 0 0 42 70
<< metal1 >>
rect 0 65 42 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 42 65
rect 0 58 42 63
rect 6 55 10 58
rect 26 55 30 58
rect 18 55 22 56
rect 6 53 7 55
rect 9 53 10 55
rect 18 53 19 55
rect 21 53 22 55
rect 26 53 27 55
rect 29 53 30 55
rect 6 51 10 53
rect 18 51 22 53
rect 26 51 30 53
rect 6 49 7 51
rect 9 49 10 51
rect 18 49 19 51
rect 21 49 22 51
rect 26 49 27 51
rect 29 49 30 51
rect 6 48 10 49
rect 18 48 22 49
rect 26 48 30 49
rect 19 46 22 48
rect 19 43 39 46
rect 36 34 39 43
rect 7 40 12 41
rect 15 40 19 41
rect 29 40 33 41
rect 7 38 8 40
rect 10 38 12 40
rect 15 38 16 40
rect 18 38 19 40
rect 29 38 30 40
rect 32 38 33 40
rect 7 37 12 38
rect 15 37 19 38
rect 29 37 33 38
rect 36 30 40 34
rect 36 19 39 30
rect 7 21 25 24
rect 7 19 10 21
rect 22 19 25 21
rect 6 18 10 19
rect 14 18 18 19
rect 22 18 26 19
rect 30 18 39 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 30 16 31 18
rect 33 16 39 18
rect 6 15 10 16
rect 14 13 18 16
rect 22 15 26 16
rect 30 15 34 16
rect 0 7 42 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 42 7
rect 0 2 42 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 7 53 9 55
rect 19 53 21 55
rect 27 53 29 55
rect 7 49 9 51
rect 19 49 21 51
rect 27 49 29 51
rect 8 38 10 40
rect 16 38 18 40
rect 30 38 32 40
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 31 16 33 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
<< poly >>
rect 11 46 13 59
rect 15 42 17 59
rect 23 42 25 59
rect 10 44 13 46
rect 10 42 12 44
rect 6 36 12 42
rect 14 38 20 42
rect 23 40 34 42
rect 27 36 34 40
rect 14 36 21 38
rect 10 27 12 36
rect 19 12 21 36
rect 27 12 29 36
rect 10 25 13 27
rect 11 12 13 25
<< ndiff >>
rect 3 61 39 67
rect 5 14 35 20
<< pdiff >>
rect 5 47 31 57
rect 3 3 39 9
<< nwell >>
rect 0 31 42 70
<< pwell >>
rect 0 0 42 31
<< end >>
