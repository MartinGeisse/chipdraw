magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577735692896
<< sizer >>
rect 0 0 49 70
<< metal1 >>
rect 0 65 49 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 49 65
rect 0 58 49 63
rect 14 55 18 58
rect 30 55 34 58
rect 6 55 10 56
rect 22 55 26 56
rect 38 55 42 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 22 53 23 55
rect 25 53 26 55
rect 30 53 31 55
rect 33 53 34 55
rect 38 53 39 55
rect 41 53 42 55
rect 6 51 10 53
rect 14 51 18 53
rect 22 51 26 53
rect 30 51 34 53
rect 38 51 42 53
rect 6 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 22 49 23 51
rect 25 49 26 51
rect 30 49 31 51
rect 33 49 34 51
rect 38 49 39 51
rect 41 49 46 51
rect 6 48 10 49
rect 14 48 18 49
rect 22 48 26 49
rect 30 48 34 49
rect 38 48 46 49
rect 7 46 10 48
rect 22 46 25 48
rect 43 41 46 48
rect 7 43 25 46
rect 15 40 18 43
rect 43 36 47 41
rect 15 39 39 40
rect 15 37 36 39
rect 38 37 39 39
rect 15 19 18 37
rect 35 36 39 37
rect 43 19 46 36
rect 1 33 12 34
rect 22 33 26 34
rect 1 31 9 33
rect 11 31 12 33
rect 22 31 23 33
rect 25 31 26 33
rect 1 30 5 31
rect 8 30 12 31
rect 22 30 26 31
rect 22 26 26 27
rect 20 25 26 26
rect 20 23 21 25
rect 23 23 26 25
rect 20 22 24 23
rect 6 18 18 19
rect 22 18 26 19
rect 30 18 46 19
rect 6 16 7 18
rect 9 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 30 16 31 18
rect 33 16 46 18
rect 6 15 10 16
rect 22 13 26 16
rect 30 15 34 16
rect 0 7 49 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 49 7
rect 0 2 49 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 7 53 9 55
rect 15 53 17 55
rect 23 53 25 55
rect 31 53 33 55
rect 39 53 41 55
rect 7 49 9 51
rect 15 49 17 51
rect 23 49 25 51
rect 31 49 33 51
rect 39 49 41 51
rect 36 37 38 39
rect 9 31 11 33
rect 23 31 25 33
rect 21 23 23 25
rect 7 16 9 18
rect 23 16 25 18
rect 31 16 33 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
<< poly >>
rect 11 35 13 59
rect 19 35 21 59
rect 27 41 29 59
rect 35 41 37 59
rect 27 39 31 41
rect 34 35 40 41
rect 29 27 31 39
rect 7 29 13 35
rect 19 31 27 35
rect 35 23 37 35
rect 15 29 27 31
rect 11 12 13 29
rect 15 12 17 29
rect 19 25 31 27
rect 19 21 25 25
rect 27 21 37 23
rect 19 12 21 21
rect 27 12 29 21
<< ndiff >>
rect 3 61 46 67
rect 5 14 35 20
<< pdiff >>
rect 5 47 43 57
rect 3 3 46 9
<< nwell >>
rect 0 31 49 70
<< pwell >>
rect 0 0 49 31
<< end >>
