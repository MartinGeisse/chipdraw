magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577095071989
<< sizer >>
rect 0 0 35 70
<< metal1 >>
rect 0 65 35 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 35 65
rect 0 58 35 63
rect 6 55 10 58
rect 22 55 26 58
rect 14 55 18 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 22 53 23 55
rect 25 53 26 55
rect 6 51 10 53
rect 14 51 18 53
rect 22 51 26 53
rect 6 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 22 49 23 51
rect 25 49 26 51
rect 6 47 10 49
rect 14 47 18 49
rect 22 47 26 49
rect 6 45 7 47
rect 9 45 10 47
rect 14 45 15 47
rect 17 45 18 47
rect 22 45 23 47
rect 25 45 26 47
rect 6 43 10 45
rect 14 43 18 45
rect 22 43 26 45
rect 6 41 7 43
rect 9 41 10 43
rect 14 41 15 43
rect 17 41 18 43
rect 22 41 23 43
rect 25 41 26 43
rect 6 40 10 41
rect 14 34 18 41
rect 22 40 26 41
rect 1 33 12 34
rect 14 30 19 34
rect 22 33 26 34
rect 1 31 9 33
rect 11 31 12 33
rect 22 31 23 33
rect 25 31 26 33
rect 1 30 5 31
rect 8 30 12 31
rect 22 30 26 31
rect 14 23 18 30
rect 6 22 10 23
rect 14 22 22 23
rect 6 20 7 22
rect 9 20 10 22
rect 14 20 19 22
rect 21 20 22 22
rect 6 18 10 20
rect 18 18 22 20
rect 6 16 7 18
rect 9 16 10 18
rect 18 16 19 18
rect 21 16 22 18
rect 6 13 10 16
rect 18 15 22 16
rect 0 7 35 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 35 7
rect 0 2 35 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 7 53 9 55
rect 15 53 17 55
rect 23 53 25 55
rect 7 49 9 51
rect 15 49 17 51
rect 23 49 25 51
rect 7 45 9 47
rect 15 45 17 47
rect 23 45 25 47
rect 7 41 9 43
rect 15 41 17 43
rect 23 41 25 43
rect 9 31 11 33
rect 23 31 25 33
rect 7 20 9 22
rect 19 20 21 22
rect 7 16 9 18
rect 19 16 21 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
<< poly >>
rect 11 35 13 59
rect 19 35 21 59
rect 7 29 13 35
rect 19 29 27 35
rect 11 12 13 29
rect 19 27 21 29
rect 15 25 21 27
rect 15 12 17 25
<< ndiff >>
rect 3 61 29 67
rect 5 14 23 24
<< pdiff >>
rect 5 39 27 57
rect 3 3 29 9
<< nwell >>
rect 0 31 35 70
<< pwell >>
rect 0 0 35 31
<< end >>
