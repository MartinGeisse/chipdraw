magic
tech concept
timestamp 1576567466492
<< sizer >>
rect 0 0 42 140
<< metal1 >>
rect 0 134 42 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 28 134
rect 30 132 32 134
rect 34 132 42 134
rect 0 128 42 132
rect 9 124 13 128
rect 29 90 32 128
rect 21 124 25 125
rect 9 122 10 124
rect 12 122 13 124
rect 21 122 22 124
rect 24 122 25 124
rect 9 120 13 122
rect 21 120 25 122
rect 9 118 10 120
rect 12 118 13 120
rect 21 118 22 120
rect 24 118 25 120
rect 9 117 13 118
rect 21 117 25 118
rect 22 100 25 117
rect 11 113 15 114
rect 2 111 12 113
rect 14 111 15 113
rect 2 110 15 111
rect 2 90 5 110
rect 15 105 19 106
rect 8 103 16 105
rect 18 103 19 105
rect 8 102 19 103
rect 8 76 11 102
rect 15 97 25 100
rect 15 48 18 97
rect 1 86 5 90
rect 22 87 32 90
rect 22 62 25 87
rect 2 31 5 86
rect 8 72 12 76
rect 8 36 11 72
rect 21 61 25 62
rect 29 61 33 62
rect 21 59 22 61
rect 24 59 25 61
rect 29 59 30 61
rect 32 59 33 61
rect 21 57 25 59
rect 29 57 33 59
rect 21 55 22 57
rect 24 55 25 57
rect 29 55 30 57
rect 32 55 33 57
rect 21 54 25 55
rect 29 54 33 55
rect 30 40 33 54
rect 15 47 21 48
rect 15 45 18 47
rect 20 45 21 47
rect 15 44 21 45
rect 18 25 21 44
rect 36 40 40 41
rect 29 39 40 40
rect 29 37 30 39
rect 32 37 40 39
rect 29 36 33 37
rect 8 33 14 36
rect 11 31 14 33
rect 29 31 34 32
rect 2 30 7 31
rect 11 30 15 31
rect 29 29 30 31
rect 32 29 34 31
rect 2 28 4 30
rect 6 28 7 30
rect 11 28 12 30
rect 14 28 15 30
rect 29 28 34 29
rect 2 27 7 28
rect 11 27 15 28
rect 31 13 34 28
rect 10 22 28 25
rect 10 20 13 22
rect 25 20 28 22
rect 9 19 13 20
rect 17 19 21 20
rect 25 19 29 20
rect 9 17 10 19
rect 12 17 13 19
rect 17 17 18 19
rect 20 17 21 19
rect 25 17 26 19
rect 28 17 29 19
rect 9 16 13 17
rect 17 13 21 17
rect 25 16 29 17
rect 0 8 42 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 28 8
rect 30 6 32 8
rect 34 6 42 8
rect 0 2 42 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 28 132 30 134
rect 32 132 34 134
rect 10 122 12 124
rect 22 122 24 124
rect 10 118 12 120
rect 22 118 24 120
rect 12 111 14 113
rect 16 103 18 105
rect 22 59 24 61
rect 30 59 32 61
rect 22 55 24 57
rect 30 55 32 57
rect 18 45 20 47
rect 30 37 32 39
rect 30 29 32 31
rect 4 28 6 30
rect 12 28 14 30
rect 10 17 12 19
rect 18 17 20 19
rect 26 17 28 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
rect 28 6 30 8
rect 32 6 34 8
<< poly >>
rect 14 115 16 128
rect 18 107 20 128
rect 10 109 16 115
rect 14 101 20 107
rect 26 52 28 65
rect 20 50 28 52
rect 20 49 22 50
rect 16 43 22 49
rect 20 35 22 43
rect 20 33 36 35
rect 2 26 8 32
rect 10 28 16 32
rect 10 26 20 28
rect 2 24 4 26
rect 18 24 20 26
rect 2 22 16 24
rect 18 22 24 24
rect 14 13 16 22
rect 22 13 24 22
<< ndiff >>
rect 6 130 36 136
rect 28 27 34 41
rect 8 15 30 21
<< pdiff >>
rect 8 116 28 126
rect 20 53 34 63
rect 6 4 36 10
<< nwell >>
rect 3 48 39 139
<< pwell >>
rect 3 1 39 46
<< end >>
