magic
tech concept
timestamp 1576404084682
<< sizer >>
rect 0 0 48 140
<< metal1 >>
rect 10 134 48 139
rect 10 132 17 134
rect 19 132 22 134
rect 24 132 27 134
rect 29 132 48 134
rect 10 128 48 132
rect 18 124 22 128
rect 26 124 30 125
rect 18 122 19 124
rect 21 122 22 124
rect 26 122 27 124
rect 29 122 30 124
rect 18 120 22 122
rect 26 120 30 122
rect 18 118 19 120
rect 21 118 22 120
rect 26 118 27 120
rect 29 118 30 120
rect 18 116 22 118
rect 26 116 30 118
rect 18 114 19 116
rect 21 114 22 116
rect 26 114 27 116
rect 29 114 30 116
rect 18 112 22 114
rect 26 112 30 114
rect 18 110 19 112
rect 21 110 22 112
rect 26 110 27 112
rect 29 110 30 112
rect 18 108 22 110
rect 26 108 30 110
rect 18 106 19 108
rect 21 106 22 108
rect 26 106 27 108
rect 29 106 30 108
rect 18 104 22 106
rect 26 104 30 106
rect 18 102 19 104
rect 21 102 22 104
rect 26 102 27 104
rect 29 102 30 104
rect 18 100 22 102
rect 26 100 30 102
rect 18 98 19 100
rect 21 98 22 100
rect 26 98 27 100
rect 29 98 30 100
rect 18 96 22 98
rect 26 96 30 98
rect 18 94 19 96
rect 21 94 22 96
rect 26 94 27 96
rect 29 94 30 96
rect 18 93 22 94
rect 26 76 30 94
rect 18 67 22 76
rect 26 72 36 76
rect 26 31 30 72
rect 18 65 19 67
rect 21 65 22 67
rect 18 64 22 65
rect 18 31 22 32
rect 18 29 19 31
rect 21 29 22 31
rect 26 29 27 31
rect 29 29 30 31
rect 18 27 22 29
rect 26 27 30 29
rect 18 25 19 27
rect 21 25 22 27
rect 26 25 27 27
rect 29 25 30 27
rect 18 23 22 25
rect 26 23 30 25
rect 18 21 19 23
rect 21 21 22 23
rect 26 21 27 23
rect 29 21 30 23
rect 18 19 22 21
rect 26 19 30 21
rect 18 17 19 19
rect 21 17 22 19
rect 26 17 27 19
rect 29 17 30 19
rect 18 13 22 17
rect 26 16 30 17
rect 10 8 38 13
rect 10 6 17 8
rect 19 6 22 8
rect 24 6 27 8
rect 29 6 38 8
rect 10 2 38 6
<< contact >>
rect 17 132 19 134
rect 22 132 24 134
rect 27 132 29 134
rect 19 122 21 124
rect 27 122 29 124
rect 19 118 21 120
rect 27 118 29 120
rect 19 114 21 116
rect 27 114 29 116
rect 19 110 21 112
rect 27 110 29 112
rect 19 106 21 108
rect 27 106 29 108
rect 19 102 21 104
rect 27 102 29 104
rect 19 98 21 100
rect 27 98 29 100
rect 19 94 21 96
rect 27 94 29 96
rect 19 65 21 67
rect 19 29 21 31
rect 27 29 29 31
rect 19 25 21 27
rect 27 25 29 27
rect 19 21 21 23
rect 27 21 29 23
rect 19 17 21 19
rect 27 17 29 19
rect 17 6 19 8
rect 22 6 24 8
rect 27 6 29 8
<< poly >>
rect 23 69 25 128
rect 17 63 25 69
rect 23 13 25 63
<< ndiff >>
rect 15 130 33 136
rect 17 15 31 33
<< pdiff >>
rect 17 92 31 126
rect 15 4 33 10
<< nwell >>
rect 12 48 36 139
<< pwell >>
rect 12 1 36 46
<< end >>
