magic
tech concept
timestamp 1576565593541
<< sizer >>
rect 0 0 42 140
<< metal1 >>
rect 0 134 42 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 28 134
rect 30 132 32 134
rect 34 132 42 134
rect 0 128 42 132
rect 11 124 15 128
rect 23 124 28 125
rect 11 122 12 124
rect 14 122 15 124
rect 23 122 24 124
rect 26 122 28 124
rect 11 120 15 122
rect 23 121 28 122
rect 23 120 30 121
rect 11 118 12 120
rect 14 118 15 120
rect 23 118 24 120
rect 26 118 30 120
rect 11 117 15 118
rect 23 117 30 118
rect 27 76 30 117
rect 13 105 17 106
rect 9 103 14 105
rect 16 103 17 105
rect 9 102 17 103
rect 9 90 12 102
rect 8 86 12 90
rect 9 36 12 86
rect 27 69 33 76
rect 30 25 33 69
rect 15 61 25 62
rect 15 59 22 61
rect 24 59 25 61
rect 15 58 25 59
rect 9 35 19 36
rect 9 33 16 35
rect 18 33 19 35
rect 15 32 19 33
rect 13 22 33 25
rect 13 19 17 22
rect 29 19 33 22
rect 21 19 25 20
rect 13 17 14 19
rect 16 17 17 19
rect 21 17 22 19
rect 24 17 25 19
rect 29 17 30 19
rect 32 17 33 19
rect 13 16 17 17
rect 21 13 25 17
rect 29 16 33 17
rect 0 8 42 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 28 8
rect 30 6 32 8
rect 34 6 42 8
rect 0 2 42 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 28 132 30 134
rect 32 132 34 134
rect 12 122 14 124
rect 24 122 26 124
rect 12 118 14 120
rect 24 118 26 120
rect 14 103 16 105
rect 22 59 24 61
rect 16 33 18 35
rect 14 17 16 19
rect 22 17 24 19
rect 30 17 32 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
rect 28 6 30 8
rect 32 6 34 8
<< poly >>
rect 16 107 18 128
rect 20 63 22 128
rect 12 101 18 107
rect 20 57 28 63
rect 26 13 28 57
rect 14 31 20 37
rect 18 13 20 31
<< ndiff >>
rect 6 130 36 136
rect 12 15 34 21
<< pdiff >>
rect 10 116 28 126
rect 6 4 36 10
<< nwell >>
rect 3 48 39 139
<< pwell >>
rect 3 1 39 46
<< end >>
