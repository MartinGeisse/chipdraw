magic
tech concept
timestamp 1576424329639
<< sizer >>
rect 0 0 42 140
<< metal1 >>
rect 0 134 42 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 28 134
rect 30 132 32 134
rect 34 132 42 134
rect 0 128 42 132
rect 19 124 23 128
rect 10 124 14 125
rect 28 124 32 125
rect 10 122 11 124
rect 13 122 14 124
rect 19 122 20 124
rect 22 122 23 124
rect 28 122 29 124
rect 31 122 32 124
rect 10 120 14 122
rect 19 120 23 122
rect 28 120 32 122
rect 10 118 11 120
rect 13 118 14 120
rect 19 118 20 120
rect 22 118 23 120
rect 28 118 29 120
rect 31 118 32 120
rect 10 117 14 118
rect 19 117 23 118
rect 28 76 32 118
rect 11 114 14 117
rect 11 113 26 114
rect 11 111 23 113
rect 25 111 26 113
rect 22 110 26 111
rect 23 27 26 110
rect 8 75 17 76
rect 28 72 33 76
rect 8 73 14 75
rect 16 73 17 75
rect 8 72 17 73
rect 28 19 32 72
rect 22 26 26 27
rect 11 24 23 26
rect 25 24 26 26
rect 11 23 26 24
rect 11 20 14 23
rect 10 19 14 20
rect 19 19 23 20
rect 10 17 11 19
rect 13 17 14 19
rect 19 17 20 19
rect 22 17 23 19
rect 28 17 29 19
rect 31 17 32 19
rect 10 16 14 17
rect 19 13 23 17
rect 28 16 32 17
rect 0 8 42 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 28 8
rect 30 6 32 8
rect 34 6 42 8
rect 0 2 42 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 28 132 30 134
rect 32 132 34 134
rect 11 122 13 124
rect 20 122 22 124
rect 29 122 31 124
rect 11 118 13 120
rect 20 118 22 120
rect 29 118 31 120
rect 23 111 25 113
rect 14 73 16 75
rect 23 24 25 26
rect 11 17 13 19
rect 20 17 22 19
rect 29 17 31 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
rect 28 6 30 8
rect 32 6 34 8
<< poly >>
rect 15 77 17 128
rect 25 115 27 128
rect 21 109 27 115
rect 12 71 18 77
rect 15 13 17 71
rect 21 22 27 28
rect 25 13 27 22
<< ndiff >>
rect 6 130 36 136
rect 9 15 33 21
<< pdiff >>
rect 9 116 33 126
rect 6 4 36 10
<< nwell >>
rect 3 48 39 139
<< pwell >>
rect 3 1 39 46
<< end >>
