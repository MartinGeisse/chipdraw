magic
tech concept
timestamp 1576654645161
<< sizer >>
rect 0 0 42 140
<< metal1 >>
rect 0 134 42 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 28 134
rect 30 132 32 134
rect 34 132 42 134
rect 0 128 42 132
rect 13 124 17 128
rect 25 124 30 125
rect 13 122 14 124
rect 16 122 17 124
rect 25 122 26 124
rect 28 122 30 124
rect 13 120 17 122
rect 25 120 30 122
rect 13 118 14 120
rect 16 118 17 120
rect 25 118 26 120
rect 28 118 30 120
rect 13 117 17 118
rect 25 117 30 118
rect 27 76 30 117
rect 15 111 19 112
rect 9 109 16 111
rect 18 109 19 111
rect 9 108 19 109
rect 9 90 12 108
rect 15 103 19 104
rect 15 102 25 103
rect 15 100 22 102
rect 24 100 25 102
rect 21 99 25 100
rect 8 86 12 90
rect 9 29 12 86
rect 27 72 33 76
rect 27 20 30 72
rect 15 40 25 41
rect 15 38 22 40
rect 24 38 25 40
rect 15 37 25 38
rect 9 28 19 29
rect 9 26 16 28
rect 18 26 19 28
rect 9 25 19 26
rect 13 19 17 20
rect 25 19 30 20
rect 13 17 14 19
rect 16 17 17 19
rect 25 17 26 19
rect 28 17 30 19
rect 13 13 17 17
rect 25 16 30 17
rect 0 8 42 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 28 8
rect 30 6 32 8
rect 34 6 42 8
rect 0 2 42 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 28 132 30 134
rect 32 132 34 134
rect 14 122 16 124
rect 26 122 28 124
rect 14 118 16 120
rect 26 118 28 120
rect 16 109 18 111
rect 22 100 24 102
rect 22 38 24 40
rect 16 26 18 28
rect 14 17 16 19
rect 26 17 28 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
rect 28 6 30 8
rect 32 6 34 8
<< poly >>
rect 18 113 20 128
rect 22 104 24 128
rect 13 106 20 113
rect 20 98 26 104
rect 20 36 26 42
rect 22 13 24 36
rect 14 24 20 30
rect 18 13 20 24
<< ndiff >>
rect 6 130 36 136
rect 12 15 30 21
<< pdiff >>
rect 12 116 30 126
rect 6 4 36 10
<< nwell >>
rect 3 48 39 139
<< pwell >>
rect 3 1 39 46
<< end >>
