magic
tech concept
timestamp 1577180690223
<< sizer >>
rect 0 0 49 70
<< metal1 >>
rect 0 65 49 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 49 65
rect 0 58 49 63
rect 6 55 10 58
rect 22 55 31 58
rect 14 55 18 56
rect 35 55 39 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 22 53 23 55
rect 25 53 28 55
rect 30 53 31 55
rect 35 53 36 55
rect 38 53 39 55
rect 6 51 10 53
rect 14 51 18 53
rect 22 51 31 53
rect 35 51 39 53
rect 6 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 22 49 23 51
rect 25 49 28 51
rect 30 49 31 51
rect 35 49 36 51
rect 38 49 39 51
rect 6 48 10 49
rect 14 46 18 49
rect 22 48 31 49
rect 35 34 39 49
rect 14 43 22 46
rect 19 35 22 43
rect 8 40 14 41
rect 8 38 11 40
rect 13 38 14 40
rect 8 37 14 38
rect 19 34 33 35
rect 1 33 6 34
rect 19 32 30 34
rect 32 32 33 34
rect 35 30 40 34
rect 1 31 3 33
rect 5 31 6 33
rect 19 23 22 32
rect 29 31 33 32
rect 1 30 6 31
rect 35 18 39 30
rect 18 18 22 23
rect 6 18 10 19
rect 27 18 31 19
rect 6 16 7 18
rect 9 16 10 18
rect 18 16 19 18
rect 21 16 22 18
rect 27 16 28 18
rect 30 16 31 18
rect 35 16 36 18
rect 38 16 39 18
rect 6 13 10 16
rect 18 15 22 16
rect 27 13 31 16
rect 35 15 39 16
rect 0 7 49 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 49 7
rect 0 2 49 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 7 53 9 55
rect 15 53 17 55
rect 23 53 25 55
rect 28 53 30 55
rect 36 53 38 55
rect 7 49 9 51
rect 15 49 17 51
rect 23 49 25 51
rect 28 49 30 51
rect 36 49 38 51
rect 11 38 13 40
rect 30 32 32 34
rect 3 31 5 33
rect 7 16 9 18
rect 19 16 21 18
rect 28 16 30 18
rect 36 16 38 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
<< poly >>
rect 11 46 13 59
rect 19 46 21 59
rect 32 36 34 59
rect 1 44 13 46
rect 15 44 21 46
rect 1 35 3 44
rect 15 42 17 44
rect 9 40 17 42
rect 9 36 15 40
rect 13 27 15 36
rect 28 30 34 36
rect 1 29 7 35
rect 32 12 34 30
rect 1 23 3 29
rect 13 25 17 27
rect 15 12 17 25
rect 1 21 13 23
rect 11 12 13 21
<< ndiff >>
rect 3 61 45 67
rect 5 14 23 20
rect 26 14 40 20
<< pdiff >>
rect 5 47 40 57
rect 3 3 45 9
<< nwell >>
rect 0 31 49 70
rect 20 29 49 31
<< pwell >>
rect 0 29 20 31
rect 0 0 49 29
<< end >>
