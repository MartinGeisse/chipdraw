magic
tech concept
timestamp 1577105533279
<< sizer >>
rect 0 0 45 70
<< metal1 >>
rect 0 65 45 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 45 65
rect 0 58 45 63
rect 6 55 10 58
rect 18 55 22 56
rect 27 55 31 56
rect 35 55 39 56
rect 6 53 7 55
rect 9 53 10 55
rect 18 53 19 55
rect 21 53 22 55
rect 27 53 28 55
rect 30 53 31 55
rect 35 53 36 55
rect 38 53 39 55
rect 6 51 10 53
rect 18 51 22 53
rect 27 51 31 53
rect 35 51 39 53
rect 6 49 7 51
rect 9 49 10 51
rect 18 49 19 51
rect 21 49 22 51
rect 27 49 28 51
rect 30 49 31 51
rect 35 49 36 51
rect 38 49 39 51
rect 6 48 10 49
rect 18 48 22 49
rect 27 47 31 49
rect 35 47 39 49
rect 19 36 22 48
rect 27 45 28 47
rect 30 45 31 47
rect 35 45 36 47
rect 38 45 39 47
rect 27 43 31 45
rect 35 43 39 45
rect 27 41 28 43
rect 30 41 31 43
rect 35 41 36 43
rect 38 41 39 43
rect 8 40 14 41
rect 27 40 31 41
rect 35 34 39 41
rect 8 38 11 40
rect 13 38 14 40
rect 8 37 14 38
rect 19 35 28 36
rect 19 33 25 35
rect 27 33 28 35
rect 1 33 6 34
rect 35 30 40 34
rect 1 31 3 33
rect 5 31 6 33
rect 19 32 28 33
rect 19 24 22 32
rect 1 30 6 31
rect 35 28 39 30
rect 31 27 39 28
rect 31 25 32 27
rect 34 25 36 27
rect 38 25 39 27
rect 31 24 39 25
rect 14 21 22 24
rect 14 18 18 21
rect 31 19 39 20
rect 6 18 10 19
rect 22 18 26 19
rect 31 17 32 19
rect 34 17 36 19
rect 38 17 39 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 31 16 39 17
rect 6 13 10 16
rect 14 15 18 16
rect 22 13 26 16
rect 0 7 45 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 45 7
rect 0 2 45 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 7 53 9 55
rect 19 53 21 55
rect 28 53 30 55
rect 36 53 38 55
rect 7 49 9 51
rect 19 49 21 51
rect 28 49 30 51
rect 36 49 38 51
rect 28 45 30 47
rect 36 45 38 47
rect 28 41 30 43
rect 36 41 38 43
rect 11 38 13 40
rect 25 33 27 35
rect 3 31 5 33
rect 32 25 34 27
rect 36 25 38 27
rect 32 17 34 19
rect 36 17 38 19
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
<< poly >>
rect 11 46 13 59
rect 15 42 17 59
rect 32 37 34 59
rect 4 44 13 46
rect 4 35 6 44
rect 9 36 17 42
rect 23 35 34 37
rect 15 23 17 36
rect 1 29 7 35
rect 23 31 29 35
rect 27 23 29 31
rect 4 23 6 29
rect 4 21 13 23
rect 15 21 21 23
rect 27 21 42 23
rect 11 12 13 21
rect 19 12 21 21
<< ndiff >>
rect 3 61 41 67
rect 30 15 40 29
rect 5 14 27 20
<< pdiff >>
rect 5 47 23 57
rect 26 39 40 57
rect 3 3 41 9
<< nwell >>
rect 0 34 45 70
rect 0 31 25 34
<< pwell >>
rect 25 31 45 34
rect 0 0 45 31
<< end >>
