magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577817382847
<< sizer >>
rect 0 0 77 70
<< metal1 >>
rect 0 65 77 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 45 65
rect 47 63 49 65
rect 51 63 53 65
rect 55 63 57 65
rect 59 63 61 65
rect 63 63 65 65
rect 67 63 69 65
rect 71 63 77 65
rect 0 58 77 63
rect 14 50 18 58
rect 42 50 46 58
rect 50 53 70 56
rect 50 50 54 53
rect 66 50 70 53
rect 6 50 10 51
rect 22 50 26 51
rect 34 50 38 51
rect 58 50 62 51
rect 6 48 7 50
rect 9 48 10 50
rect 14 48 15 50
rect 17 48 18 50
rect 22 48 23 50
rect 25 48 26 50
rect 34 48 35 50
rect 37 48 38 50
rect 42 48 43 50
rect 45 48 46 50
rect 50 48 51 50
rect 53 48 54 50
rect 58 48 59 50
rect 61 48 62 50
rect 66 48 67 50
rect 69 48 70 50
rect 6 46 10 48
rect 14 46 18 48
rect 22 47 26 48
rect 34 46 38 48
rect 42 46 46 48
rect 50 46 54 48
rect 58 46 62 48
rect 66 46 70 48
rect 22 46 31 47
rect 1 44 7 46
rect 9 44 10 46
rect 14 44 15 46
rect 17 44 18 46
rect 22 44 23 46
rect 25 44 31 46
rect 34 44 35 46
rect 37 44 38 46
rect 42 44 43 46
rect 45 44 46 46
rect 50 44 51 46
rect 53 44 54 46
rect 58 44 59 46
rect 61 44 62 46
rect 66 44 67 46
rect 69 44 70 46
rect 1 43 10 44
rect 14 43 18 44
rect 22 43 31 44
rect 34 41 38 44
rect 42 43 46 44
rect 50 41 54 44
rect 58 43 62 44
rect 66 43 70 44
rect 1 28 4 43
rect 28 36 31 43
rect 59 41 62 43
rect 34 38 54 41
rect 59 38 74 41
rect 71 34 74 38
rect 28 34 67 36
rect 8 33 12 34
rect 15 33 20 34
rect 28 33 68 34
rect 71 30 75 34
rect 8 31 9 33
rect 11 31 12 33
rect 15 31 17 33
rect 19 31 20 33
rect 64 31 65 33
rect 67 31 68 33
rect 8 30 12 31
rect 15 30 20 31
rect 23 30 52 31
rect 64 30 68 31
rect 23 28 49 30
rect 51 28 52 30
rect 64 29 67 30
rect 71 24 74 30
rect 55 26 67 29
rect 1 25 26 28
rect 48 27 52 28
rect 55 24 58 26
rect 1 19 4 25
rect 37 21 58 24
rect 61 21 74 24
rect 37 19 40 21
rect 61 19 64 21
rect 1 18 10 19
rect 14 18 18 19
rect 22 18 40 19
rect 42 18 46 19
rect 54 18 64 19
rect 66 18 70 19
rect 1 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 40 18
rect 42 16 43 18
rect 45 16 46 18
rect 54 16 55 18
rect 57 16 64 18
rect 66 16 67 18
rect 69 16 70 18
rect 6 15 10 16
rect 14 13 18 16
rect 22 15 26 16
rect 42 13 46 16
rect 54 15 58 16
rect 66 13 70 16
rect 0 7 77 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 45 7
rect 47 5 49 7
rect 51 5 53 7
rect 55 5 57 7
rect 59 5 61 7
rect 63 5 65 7
rect 67 5 69 7
rect 71 5 77 7
rect 0 2 77 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 45 63 47 65
rect 49 63 51 65
rect 53 63 55 65
rect 57 63 59 65
rect 61 63 63 65
rect 65 63 67 65
rect 69 63 71 65
rect 7 48 9 50
rect 15 48 17 50
rect 23 48 25 50
rect 35 48 37 50
rect 43 48 45 50
rect 51 48 53 50
rect 59 48 61 50
rect 67 48 69 50
rect 7 44 9 46
rect 15 44 17 46
rect 23 44 25 46
rect 35 44 37 46
rect 43 44 45 46
rect 51 44 53 46
rect 59 44 61 46
rect 67 44 69 46
rect 9 31 11 33
rect 17 31 19 33
rect 65 31 67 33
rect 49 28 51 30
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 43 16 45 18
rect 55 16 57 18
rect 67 16 69 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
rect 45 5 47 7
rect 49 5 51 7
rect 53 5 55 7
rect 57 5 59 7
rect 61 5 63 7
rect 65 5 67 7
rect 69 5 71 7
<< poly >>
rect 11 56 57 58
rect 11 35 13 56
rect 55 41 57 56
rect 19 35 21 54
rect 39 33 41 54
rect 47 32 49 54
rect 63 35 65 54
rect 55 39 61 41
rect 59 12 61 39
rect 7 29 13 35
rect 15 33 21 35
rect 63 29 70 35
rect 15 31 41 33
rect 47 26 53 32
rect 15 29 21 31
rect 39 23 41 31
rect 11 12 13 29
rect 19 12 21 29
rect 63 12 65 29
rect 51 12 53 26
rect 39 21 49 23
rect 47 12 49 21
<< ndiff >>
rect 3 61 74 67
rect 5 14 27 20
rect 41 14 71 20
<< pdiff >>
rect 5 42 27 52
rect 33 42 71 52
rect 3 3 74 9
<< nwell >>
rect 0 31 77 70
<< pwell >>
rect 0 0 77 31
<< end >>
