magic
tech concept
timestamp 1577260060035
<< sizer >>
rect 0 0 49 70
<< metal1 >>
rect 0 65 49 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 49 65
rect 0 58 49 63
rect 6 55 10 58
rect 22 55 26 58
rect 38 55 42 58
rect 14 55 18 56
rect 30 55 34 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 22 53 23 55
rect 25 53 26 55
rect 30 53 31 55
rect 33 53 34 55
rect 38 53 39 55
rect 41 53 42 55
rect 6 51 10 53
rect 14 51 18 53
rect 22 51 26 53
rect 30 51 34 53
rect 38 51 42 53
rect 6 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 22 49 23 51
rect 25 49 26 51
rect 30 49 31 51
rect 33 49 34 51
rect 38 49 39 51
rect 41 49 42 51
rect 6 48 10 49
rect 14 46 18 49
rect 22 48 26 49
rect 30 46 34 49
rect 38 48 42 49
rect 14 43 42 46
rect 39 41 42 43
rect 15 40 20 41
rect 22 40 28 41
rect 39 37 47 41
rect 15 38 17 40
rect 19 38 20 40
rect 22 38 25 40
rect 27 38 28 40
rect 15 37 20 38
rect 22 37 28 38
rect 39 18 42 37
rect 1 33 12 34
rect 28 32 33 34
rect 1 31 9 33
rect 11 31 12 33
rect 28 30 29 32
rect 31 30 33 32
rect 1 30 5 31
rect 8 30 12 31
rect 28 29 33 30
rect 6 22 10 23
rect 26 22 30 23
rect 6 20 7 22
rect 9 20 10 22
rect 26 20 27 22
rect 29 20 30 22
rect 6 18 10 20
rect 26 18 30 20
rect 6 16 7 18
rect 9 16 10 18
rect 26 16 27 18
rect 29 16 42 18
rect 6 13 10 16
rect 26 15 42 16
rect 0 7 49 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 49 7
rect 0 2 49 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 7 53 9 55
rect 15 53 17 55
rect 23 53 25 55
rect 31 53 33 55
rect 39 53 41 55
rect 7 49 9 51
rect 15 49 17 51
rect 23 49 25 51
rect 31 49 33 51
rect 39 49 41 51
rect 17 38 19 40
rect 25 38 27 40
rect 9 31 11 33
rect 29 30 31 32
rect 7 20 9 22
rect 27 20 29 22
rect 7 16 9 18
rect 27 16 29 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
<< poly >>
rect 11 35 13 59
rect 19 42 21 59
rect 27 42 29 59
rect 35 45 37 59
rect 31 43 37 45
rect 31 34 33 43
rect 15 36 21 42
rect 23 36 29 42
rect 15 12 17 36
rect 23 34 25 36
rect 7 29 13 35
rect 19 32 25 34
rect 27 30 33 34
rect 19 12 21 32
rect 23 28 33 30
rect 11 12 13 29
rect 23 12 25 28
<< ndiff >>
rect 3 61 45 67
rect 5 14 31 24
<< pdiff >>
rect 5 47 43 57
rect 3 3 45 9
<< nwell >>
rect 0 31 49 70
<< pwell >>
rect 0 0 49 31
<< end >>
