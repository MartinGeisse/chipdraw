magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577182806882
<< sizer >>
rect 0 0 49 70
<< metal1 >>
rect 0 65 49 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 49 65
rect 0 58 49 63
rect 6 55 10 58
rect 32 50 36 58
rect 18 55 22 56
rect 6 53 7 55
rect 9 53 10 55
rect 18 53 19 55
rect 21 53 22 55
rect 6 51 10 53
rect 18 51 22 53
rect 6 49 7 51
rect 9 49 10 51
rect 18 49 19 51
rect 21 49 22 51
rect 32 48 33 50
rect 35 48 36 50
rect 6 48 10 49
rect 18 48 22 49
rect 19 36 22 48
rect 32 47 36 48
rect 32 42 36 43
rect 32 40 33 42
rect 35 40 36 42
rect 8 40 14 41
rect 8 38 11 40
rect 13 38 14 40
rect 32 34 36 40
rect 8 37 14 38
rect 19 35 29 36
rect 19 33 26 35
rect 28 33 29 35
rect 1 33 6 34
rect 32 30 41 34
rect 1 31 3 33
rect 5 31 6 33
rect 19 32 29 33
rect 19 24 22 32
rect 1 30 6 31
rect 32 26 36 30
rect 32 24 33 26
rect 35 24 36 26
rect 14 21 22 24
rect 32 23 36 24
rect 14 18 18 21
rect 6 18 10 19
rect 22 18 26 19
rect 32 18 36 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 32 16 33 18
rect 35 16 36 18
rect 6 13 10 16
rect 14 15 18 16
rect 22 13 26 16
rect 32 13 36 16
rect 0 7 49 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 49 7
rect 0 2 49 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 7 53 9 55
rect 19 53 21 55
rect 7 49 9 51
rect 19 49 21 51
rect 33 48 35 50
rect 33 40 35 42
rect 11 38 13 40
rect 26 33 28 35
rect 3 31 5 33
rect 33 24 35 26
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 33 16 35 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
<< poly >>
rect 11 46 13 59
rect 15 42 17 59
rect 4 44 13 46
rect 28 44 39 46
rect 4 35 6 44
rect 28 37 30 44
rect 9 36 17 42
rect 24 31 30 37
rect 15 23 17 36
rect 1 29 7 35
rect 28 22 30 31
rect 4 23 6 29
rect 4 21 13 23
rect 15 21 21 23
rect 28 20 39 22
rect 11 12 13 21
rect 19 12 21 21
<< ndiff >>
rect 3 61 45 67
rect 31 14 37 28
rect 5 14 27 20
<< pdiff >>
rect 5 47 23 57
rect 31 38 37 52
rect 3 3 45 9
<< nwell >>
rect 0 33 49 70
rect 0 31 26 33
<< pwell >>
rect 26 31 49 33
rect 0 0 49 31
<< end >>
