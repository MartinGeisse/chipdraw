magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577171279542
<< sizer >>
rect 0 0 42 70
<< metal1 >>
rect 0 65 42 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 42 65
rect 0 58 42 63
rect 14 55 18 58
rect 6 55 10 56
rect 22 55 26 56
rect 30 55 34 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 22 53 23 55
rect 25 53 26 55
rect 30 53 31 55
rect 33 53 34 55
rect 6 51 10 53
rect 14 51 18 53
rect 22 51 26 53
rect 30 51 34 53
rect 6 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 22 49 23 51
rect 25 49 26 51
rect 30 49 31 51
rect 33 49 34 51
rect 6 46 10 49
rect 14 48 18 49
rect 22 46 26 49
rect 30 48 34 49
rect 31 32 34 48
rect 6 43 26 46
rect 8 40 12 41
rect 20 40 26 41
rect 8 38 9 40
rect 11 38 12 40
rect 20 38 21 40
rect 23 38 26 40
rect 8 37 12 38
rect 20 37 26 38
rect 19 29 34 32
rect 19 19 22 29
rect 28 26 33 27
rect 28 24 29 26
rect 31 24 33 26
rect 28 23 33 24
rect 6 18 10 19
rect 18 18 22 19
rect 26 18 30 19
rect 6 16 7 18
rect 9 16 10 18
rect 18 16 19 18
rect 21 16 22 18
rect 26 16 27 18
rect 29 16 30 18
rect 6 13 10 16
rect 18 15 22 16
rect 26 13 30 16
rect 0 7 42 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 42 7
rect 0 2 42 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 7 53 9 55
rect 15 53 17 55
rect 23 53 25 55
rect 31 53 33 55
rect 7 49 9 51
rect 15 49 17 51
rect 23 49 25 51
rect 31 49 33 51
rect 9 38 11 40
rect 21 38 23 40
rect 29 24 31 26
rect 7 16 9 18
rect 19 16 21 18
rect 27 16 29 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
<< poly >>
rect 11 42 13 59
rect 19 42 21 59
rect 27 28 29 59
rect 7 36 13 42
rect 19 36 25 42
rect 11 12 13 36
rect 19 33 21 36
rect 15 31 21 33
rect 15 12 17 31
rect 27 24 33 28
rect 23 22 33 24
rect 23 12 25 22
<< ndiff >>
rect 3 61 37 67
rect 5 14 31 20
<< pdiff >>
rect 5 47 35 57
rect 3 3 37 9
<< nwell >>
rect 0 31 42 70
<< pwell >>
rect 0 0 42 31
<< end >>
