magic
tech concept
timestamp 1576309957687
<< sizer >>
rect 0 0 28 140
<< metal1 >>
rect 0 134 28 139
rect 0 132 7 134
rect 9 132 12 134
rect 14 132 17 134
rect 19 132 28 134
rect 0 128 28 132
rect 8 124 12 128
rect 16 124 20 125
rect 8 122 9 124
rect 11 122 12 124
rect 16 122 17 124
rect 19 122 20 124
rect 8 120 12 122
rect 16 120 20 122
rect 8 118 9 120
rect 11 118 12 120
rect 16 118 17 120
rect 19 118 20 120
rect 8 116 12 118
rect 16 116 20 118
rect 8 114 9 116
rect 11 114 12 116
rect 16 114 17 116
rect 19 114 20 116
rect 8 112 12 114
rect 16 112 20 114
rect 8 110 9 112
rect 11 110 12 112
rect 16 110 17 112
rect 19 110 20 112
rect 8 108 12 110
rect 16 108 20 110
rect 8 106 9 108
rect 11 106 12 108
rect 16 106 17 108
rect 19 106 20 108
rect 8 104 12 106
rect 16 104 20 106
rect 8 102 9 104
rect 11 102 12 104
rect 16 102 17 104
rect 19 102 20 104
rect 8 100 12 102
rect 16 100 20 102
rect 8 98 9 100
rect 11 98 12 100
rect 16 98 17 100
rect 19 98 20 100
rect 8 96 12 98
rect 16 96 20 98
rect 8 94 9 96
rect 11 94 12 96
rect 16 94 17 96
rect 19 94 20 96
rect 8 93 12 94
rect 16 76 20 94
rect 8 67 12 76
rect 16 72 26 76
rect 16 31 20 72
rect 8 65 9 67
rect 11 65 12 67
rect 8 64 12 65
rect 8 31 12 32
rect 8 29 9 31
rect 11 29 12 31
rect 16 29 17 31
rect 19 29 20 31
rect 8 27 12 29
rect 16 27 20 29
rect 8 25 9 27
rect 11 25 12 27
rect 16 25 17 27
rect 19 25 20 27
rect 8 23 12 25
rect 16 23 20 25
rect 8 21 9 23
rect 11 21 12 23
rect 16 21 17 23
rect 19 21 20 23
rect 8 19 12 21
rect 16 19 20 21
rect 8 17 9 19
rect 11 17 12 19
rect 16 17 17 19
rect 19 17 20 19
rect 8 13 12 17
rect 16 16 20 17
rect 0 8 28 13
rect 0 6 7 8
rect 9 6 12 8
rect 14 6 17 8
rect 19 6 28 8
rect 0 2 28 6
<< contact >>
rect 7 132 9 134
rect 12 132 14 134
rect 17 132 19 134
rect 9 122 11 124
rect 17 122 19 124
rect 9 118 11 120
rect 17 118 19 120
rect 9 114 11 116
rect 17 114 19 116
rect 9 110 11 112
rect 17 110 19 112
rect 9 106 11 108
rect 17 106 19 108
rect 9 102 11 104
rect 17 102 19 104
rect 9 98 11 100
rect 17 98 19 100
rect 9 94 11 96
rect 17 94 19 96
rect 9 65 11 67
rect 9 29 11 31
rect 17 29 19 31
rect 9 25 11 27
rect 17 25 19 27
rect 9 21 11 23
rect 17 21 19 23
rect 9 17 11 19
rect 17 17 19 19
rect 7 6 9 8
rect 12 6 14 8
rect 17 6 19 8
<< poly >>
rect 13 69 15 128
rect 7 63 15 69
rect 13 13 15 63
<< ndiff >>
rect 5 130 23 136
rect 7 15 21 33
<< pdiff >>
rect 7 92 21 126
rect 5 4 23 10
<< nwell >>
rect 2 48 26 139
<< pwell >>
rect 2 1 26 46
<< end >>
