magic
tech concept
timestamp 1576406358155
<< sizer >>
rect 0 0 35 140
<< metal1 >>
rect 0 134 35 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 35 134
rect 0 128 35 132
rect 11 124 15 128
rect 19 124 23 125
rect 11 122 12 124
rect 14 122 15 124
rect 19 122 20 124
rect 22 122 23 124
rect 11 120 15 122
rect 19 120 23 122
rect 11 118 12 120
rect 14 118 15 120
rect 19 118 20 120
rect 22 118 23 120
rect 11 116 15 118
rect 19 116 23 118
rect 11 114 12 116
rect 14 114 15 116
rect 19 114 20 116
rect 22 114 23 116
rect 11 112 15 114
rect 19 112 23 114
rect 11 110 12 112
rect 14 110 15 112
rect 19 110 20 112
rect 22 110 23 112
rect 11 108 15 110
rect 19 108 23 110
rect 11 106 12 108
rect 14 106 15 108
rect 19 106 20 108
rect 22 106 23 108
rect 11 104 15 106
rect 19 104 23 106
rect 11 102 12 104
rect 14 102 15 104
rect 19 102 20 104
rect 22 102 23 104
rect 11 100 15 102
rect 19 100 23 102
rect 11 98 12 100
rect 14 98 15 100
rect 19 98 20 100
rect 22 98 23 100
rect 11 96 15 98
rect 19 96 23 98
rect 11 94 12 96
rect 14 94 15 96
rect 19 94 20 96
rect 22 94 23 96
rect 11 93 15 94
rect 19 76 23 94
rect 8 75 17 76
rect 19 72 26 76
rect 8 73 14 75
rect 16 73 17 75
rect 8 72 17 73
rect 19 31 23 72
rect 11 31 15 32
rect 11 29 12 31
rect 14 29 15 31
rect 19 29 20 31
rect 22 29 23 31
rect 11 27 15 29
rect 19 27 23 29
rect 11 25 12 27
rect 14 25 15 27
rect 19 25 20 27
rect 22 25 23 27
rect 11 23 15 25
rect 19 23 23 25
rect 11 21 12 23
rect 14 21 15 23
rect 19 21 20 23
rect 22 21 23 23
rect 11 19 15 21
rect 19 19 23 21
rect 11 17 12 19
rect 14 17 15 19
rect 19 17 20 19
rect 22 17 23 19
rect 11 13 15 17
rect 19 16 23 17
rect 0 8 35 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 35 8
rect 0 2 35 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 12 122 14 124
rect 20 122 22 124
rect 12 118 14 120
rect 20 118 22 120
rect 12 114 14 116
rect 20 114 22 116
rect 12 110 14 112
rect 20 110 22 112
rect 12 106 14 108
rect 20 106 22 108
rect 12 102 14 104
rect 20 102 22 104
rect 12 98 14 100
rect 20 98 22 100
rect 12 94 14 96
rect 20 94 22 96
rect 14 73 16 75
rect 12 29 14 31
rect 20 29 22 31
rect 12 25 14 27
rect 20 25 22 27
rect 12 21 14 23
rect 20 21 22 23
rect 12 17 14 19
rect 20 17 22 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
<< poly >>
rect 16 77 18 128
rect 12 71 18 77
rect 16 13 18 71
<< ndiff >>
rect 6 130 29 136
rect 10 15 24 33
<< pdiff >>
rect 10 92 24 126
rect 6 4 29 10
<< nwell >>
rect 3 48 32 139
<< pwell >>
rect 3 1 32 46
<< end >>
