magic
tech concept
timestamp 1577735397456
<< sizer >>
rect 0 0 49 70
<< metal1 >>
rect 0 65 49 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 49 65
rect 0 58 49 63
rect 22 55 26 58
rect 6 55 10 56
rect 30 55 34 56
rect 6 53 7 55
rect 9 53 10 55
rect 22 53 23 55
rect 25 53 26 55
rect 30 53 31 55
rect 33 53 34 55
rect 6 51 10 53
rect 22 51 26 53
rect 30 51 34 53
rect 6 49 7 51
rect 9 49 18 51
rect 22 49 23 51
rect 25 49 26 51
rect 30 49 31 51
rect 33 49 46 51
rect 6 48 18 49
rect 22 48 26 49
rect 30 48 46 49
rect 15 44 18 48
rect 43 34 46 48
rect 34 44 38 45
rect 15 42 35 44
rect 37 42 38 44
rect 15 41 38 42
rect 15 24 18 41
rect 1 33 12 34
rect 22 33 26 34
rect 29 33 34 34
rect 43 30 47 34
rect 1 31 9 33
rect 11 31 12 33
rect 22 31 23 33
rect 25 31 26 33
rect 29 31 31 33
rect 33 31 34 33
rect 1 30 5 31
rect 8 30 12 31
rect 22 30 26 31
rect 29 30 34 31
rect 43 19 46 30
rect 7 21 25 24
rect 7 19 10 21
rect 22 19 25 21
rect 6 18 10 19
rect 14 18 18 19
rect 22 18 26 19
rect 30 18 34 19
rect 38 18 46 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 30 16 31 18
rect 33 16 34 18
rect 38 16 39 18
rect 41 16 46 18
rect 6 15 10 16
rect 14 13 18 16
rect 22 15 26 16
rect 30 13 34 16
rect 38 15 42 16
rect 0 7 49 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 49 7
rect 0 2 49 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 7 53 9 55
rect 23 53 25 55
rect 31 53 33 55
rect 7 49 9 51
rect 23 49 25 51
rect 31 49 33 51
rect 35 42 37 44
rect 9 31 11 33
rect 23 31 25 33
rect 31 31 33 33
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 31 16 33 18
rect 39 16 41 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
<< poly >>
rect 11 35 13 59
rect 15 35 17 59
rect 19 42 21 59
rect 27 46 29 59
rect 27 44 39 46
rect 33 40 39 44
rect 19 40 31 42
rect 29 35 31 40
rect 37 27 39 40
rect 7 29 13 35
rect 15 33 27 35
rect 29 29 35 35
rect 19 29 27 33
rect 11 12 13 29
rect 19 12 21 29
rect 29 25 31 29
rect 35 25 39 27
rect 27 23 31 25
rect 35 12 37 25
rect 27 12 29 23
<< ndiff >>
rect 3 61 46 67
rect 5 14 43 20
<< pdiff >>
rect 5 47 35 57
rect 3 3 46 9
<< nwell >>
rect 0 31 49 70
<< pwell >>
rect 0 0 49 31
<< end >>
