magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577734289707
<< sizer >>
rect 0 0 49 70
<< metal1 >>
rect 0 65 49 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 49 65
rect 0 58 49 63
rect 6 55 10 58
rect 26 55 30 56
rect 6 53 7 55
rect 9 53 10 55
rect 26 53 27 55
rect 29 53 30 55
rect 6 51 10 53
rect 26 51 30 53
rect 6 49 7 51
rect 9 49 10 51
rect 26 49 27 51
rect 29 49 30 51
rect 6 47 10 49
rect 26 47 30 49
rect 6 45 7 47
rect 9 45 10 47
rect 26 45 27 47
rect 29 45 46 47
rect 6 44 10 45
rect 26 44 46 45
rect 43 34 46 44
rect 1 33 12 34
rect 15 32 20 34
rect 22 32 28 34
rect 36 33 40 34
rect 43 30 47 34
rect 1 31 9 33
rect 11 31 12 33
rect 36 31 37 33
rect 39 31 40 33
rect 15 30 17 32
rect 19 30 20 32
rect 22 30 25 32
rect 27 30 28 32
rect 1 30 5 31
rect 8 30 12 31
rect 36 30 40 31
rect 15 29 20 30
rect 24 29 28 30
rect 43 24 46 30
rect 15 21 46 24
rect 15 19 18 21
rect 30 19 33 21
rect 6 18 10 19
rect 14 18 18 19
rect 22 18 26 19
rect 30 18 34 19
rect 38 18 42 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 30 16 31 18
rect 33 16 34 18
rect 38 16 39 18
rect 41 16 42 18
rect 6 13 10 16
rect 14 15 18 16
rect 22 13 26 16
rect 30 15 34 16
rect 38 13 42 16
rect 0 7 49 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 34 7
rect 36 5 38 7
rect 40 5 42 7
rect 44 5 49 7
rect 0 2 49 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 7 53 9 55
rect 27 53 29 55
rect 7 49 9 51
rect 27 49 29 51
rect 7 45 9 47
rect 27 45 29 47
rect 9 31 11 33
rect 37 31 39 33
rect 17 30 19 32
rect 25 30 27 32
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 31 16 33 18
rect 39 16 41 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 34 5 36 7
rect 38 5 40 7
rect 42 5 44 7
<< poly >>
rect 11 35 13 59
rect 15 34 17 59
rect 19 38 21 59
rect 23 42 25 59
rect 23 40 37 42
rect 35 35 37 40
rect 19 36 25 38
rect 23 34 25 36
rect 7 29 13 35
rect 35 29 41 35
rect 15 28 21 34
rect 23 28 29 34
rect 11 12 13 29
rect 35 12 37 29
rect 19 12 21 28
rect 27 12 29 28
<< ndiff >>
rect 3 61 45 67
rect 5 14 43 20
<< pdiff >>
rect 5 43 31 57
rect 3 3 46 9
<< nwell >>
rect 0 31 49 70
<< pwell >>
rect 0 0 49 31
<< end >>
