magic
tech concept
timestamp 1577104493242
<< sizer >>
rect 0 0 35 70
<< metal1 >>
rect 0 65 35 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 35 65
rect 0 58 35 63
rect 6 55 10 58
rect 18 55 22 56
rect 6 53 7 55
rect 9 53 10 55
rect 18 53 19 55
rect 21 53 22 55
rect 6 51 10 53
rect 18 51 22 53
rect 6 49 7 51
rect 9 49 10 51
rect 18 49 19 51
rect 21 49 22 51
rect 6 47 10 49
rect 18 47 22 49
rect 6 45 7 47
rect 9 45 10 47
rect 18 45 19 47
rect 21 45 22 47
rect 6 43 10 45
rect 18 43 22 45
rect 6 41 7 43
rect 9 41 10 43
rect 15 41 19 43
rect 21 41 22 43
rect 6 40 10 41
rect 15 40 22 41
rect 15 34 18 40
rect 1 33 12 34
rect 15 30 19 34
rect 22 33 26 34
rect 1 31 9 33
rect 11 31 12 33
rect 22 31 23 33
rect 25 31 26 33
rect 1 30 5 31
rect 8 30 12 31
rect 22 30 26 31
rect 15 23 18 30
rect 6 22 10 23
rect 14 22 18 23
rect 22 22 26 23
rect 6 20 7 22
rect 9 20 10 22
rect 14 20 15 22
rect 17 20 18 22
rect 22 20 23 22
rect 25 20 26 22
rect 6 18 10 20
rect 14 18 18 20
rect 22 18 26 20
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 6 13 10 16
rect 14 15 18 16
rect 22 13 26 16
rect 0 7 35 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 35 7
rect 0 2 35 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 7 53 9 55
rect 19 53 21 55
rect 7 49 9 51
rect 19 49 21 51
rect 7 45 9 47
rect 19 45 21 47
rect 7 41 9 43
rect 19 41 21 43
rect 9 31 11 33
rect 23 31 25 33
rect 7 20 9 22
rect 15 20 17 22
rect 23 20 25 22
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
<< poly >>
rect 11 35 13 59
rect 15 35 17 59
rect 7 29 13 35
rect 15 33 27 35
rect 19 29 27 33
rect 11 12 13 29
rect 19 12 21 29
<< ndiff >>
rect 3 61 29 67
rect 5 14 27 24
<< pdiff >>
rect 5 39 23 57
rect 3 3 29 9
<< nwell >>
rect 0 31 35 70
<< pwell >>
rect 0 0 35 31
<< end >>
