magic
tech concept
timestamp 1577801575525
<< sizer >>
rect 0 0 35 70
<< metal1 >>
rect 0 65 35 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 35 65
rect 0 58 35 63
rect 14 55 18 58
rect 6 55 10 56
rect 22 55 26 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 22 53 23 55
rect 25 53 26 55
rect 6 51 10 53
rect 14 51 18 53
rect 22 51 26 53
rect 2 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 22 49 23 51
rect 25 49 32 51
rect 2 48 10 49
rect 14 48 18 49
rect 22 48 32 49
rect 2 34 5 48
rect 29 34 32 48
rect 1 29 5 34
rect 8 33 12 34
rect 22 33 26 34
rect 29 29 33 34
rect 8 31 9 33
rect 11 31 12 33
rect 22 31 23 33
rect 25 31 26 33
rect 8 30 12 31
rect 22 30 26 31
rect 2 19 5 29
rect 29 19 32 29
rect 2 18 10 19
rect 14 18 18 19
rect 22 18 32 19
rect 2 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 32 18
rect 6 15 10 16
rect 14 13 18 16
rect 22 15 26 16
rect 0 7 35 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 35 7
rect 0 2 35 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 7 53 9 55
rect 15 53 17 55
rect 23 53 25 55
rect 7 49 9 51
rect 15 49 17 51
rect 23 49 25 51
rect 9 31 11 33
rect 23 31 25 33
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
<< poly >>
rect 11 35 13 59
rect 19 35 21 59
rect 7 29 13 35
rect 19 29 27 35
rect 11 12 13 29
rect 19 12 21 29
<< ndiff >>
rect 3 61 32 67
rect 5 14 27 20
<< pdiff >>
rect 5 47 27 57
rect 3 3 32 9
<< nwell >>
rect 0 31 35 70
<< pwell >>
rect 0 0 35 31
<< end >>
