magic
tech concept
timestamp 1577733934236
<< sizer >>
rect 0 0 28 70
<< metal1 >>
rect 0 65 28 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 28 65
rect 0 58 28 63
rect 6 55 10 58
rect 14 55 18 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 6 51 10 53
rect 14 51 18 53
rect 6 49 7 51
rect 9 49 10 51
rect 14 49 15 51
rect 17 49 18 51
rect 6 48 10 49
rect 14 48 18 49
rect 14 33 17 48
rect 8 33 12 34
rect 22 30 26 34
rect 8 31 9 33
rect 11 31 17 33
rect 8 30 17 31
rect 22 19 25 30
rect 6 18 10 19
rect 14 18 25 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 25 18
rect 6 13 10 16
rect 14 15 18 16
rect 0 7 28 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 28 7
rect 0 2 28 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 7 53 9 55
rect 15 53 17 55
rect 7 49 9 51
rect 15 49 17 51
rect 9 31 11 33
rect 7 16 9 18
rect 15 16 17 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
<< poly >>
rect 11 35 13 59
rect 7 29 13 35
rect 11 12 13 29
<< ndiff >>
rect 3 61 25 67
rect 5 14 19 20
<< pdiff >>
rect 5 47 19 57
rect 3 3 25 9
<< nwell >>
rect 0 31 28 70
<< pwell >>
rect 0 0 28 31
<< end >>
