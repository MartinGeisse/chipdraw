magic
tech concept
timestamp 1576407036455
<< sizer >>
rect 0 0 42 140
<< metal1 >>
rect 0 134 42 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 28 134
rect 30 132 32 134
rect 34 132 42 134
rect 0 128 42 132
rect 9 124 13 128
rect 25 124 29 128
rect 17 124 21 125
rect 9 122 10 124
rect 12 122 13 124
rect 17 122 18 124
rect 20 122 21 124
rect 25 122 26 124
rect 28 122 29 124
rect 9 120 13 122
rect 17 120 21 122
rect 25 120 29 122
rect 9 118 10 120
rect 12 118 13 120
rect 17 118 18 120
rect 20 118 21 120
rect 25 118 26 120
rect 28 118 29 120
rect 9 116 13 118
rect 17 116 21 118
rect 25 116 29 118
rect 9 114 10 116
rect 12 114 13 116
rect 17 114 18 116
rect 20 114 21 116
rect 25 114 26 116
rect 28 114 29 116
rect 9 112 13 114
rect 17 112 21 114
rect 25 112 29 114
rect 9 110 10 112
rect 12 110 13 112
rect 17 110 18 112
rect 20 110 21 112
rect 25 110 26 112
rect 28 110 29 112
rect 9 108 13 110
rect 17 108 21 110
rect 25 108 29 110
rect 9 106 10 108
rect 12 106 13 108
rect 17 106 18 108
rect 20 106 21 108
rect 25 106 26 108
rect 28 106 29 108
rect 9 104 13 106
rect 17 104 21 106
rect 25 104 29 106
rect 9 102 10 104
rect 12 102 13 104
rect 17 102 18 104
rect 20 102 21 104
rect 25 102 26 104
rect 28 102 29 104
rect 9 100 13 102
rect 17 100 21 102
rect 25 100 29 102
rect 9 98 10 100
rect 12 98 13 100
rect 17 98 18 100
rect 20 98 21 100
rect 25 98 26 100
rect 28 98 29 100
rect 9 96 13 98
rect 17 96 21 98
rect 25 96 29 98
rect 9 94 10 96
rect 12 94 13 96
rect 17 94 18 96
rect 20 94 21 96
rect 25 94 26 96
rect 28 94 29 96
rect 9 93 13 94
rect 17 83 21 94
rect 25 93 29 94
rect 17 79 25 83
rect 21 76 25 79
rect 8 75 18 76
rect 21 72 26 76
rect 8 73 14 75
rect 16 73 18 75
rect 8 72 18 73
rect 21 69 25 72
rect 17 65 25 69
rect 17 31 21 65
rect 9 31 13 32
rect 25 31 29 32
rect 9 29 10 31
rect 12 29 13 31
rect 17 29 18 31
rect 20 29 21 31
rect 25 29 26 31
rect 28 29 29 31
rect 9 27 13 29
rect 17 27 21 29
rect 25 27 29 29
rect 9 25 10 27
rect 12 25 13 27
rect 17 25 18 27
rect 20 25 21 27
rect 25 25 26 27
rect 28 25 29 27
rect 9 23 13 25
rect 17 23 21 25
rect 25 23 29 25
rect 9 21 10 23
rect 12 21 13 23
rect 17 21 18 23
rect 20 21 21 23
rect 25 21 26 23
rect 28 21 29 23
rect 9 19 13 21
rect 17 19 21 21
rect 25 19 29 21
rect 9 17 10 19
rect 12 17 13 19
rect 17 17 18 19
rect 20 17 21 19
rect 25 17 26 19
rect 28 17 29 19
rect 9 13 13 17
rect 17 16 21 17
rect 25 13 29 17
rect 0 8 42 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 28 8
rect 30 6 32 8
rect 34 6 42 8
rect 0 2 42 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 28 132 30 134
rect 32 132 34 134
rect 10 122 12 124
rect 18 122 20 124
rect 26 122 28 124
rect 10 118 12 120
rect 18 118 20 120
rect 26 118 28 120
rect 10 114 12 116
rect 18 114 20 116
rect 26 114 28 116
rect 10 110 12 112
rect 18 110 20 112
rect 26 110 28 112
rect 10 106 12 108
rect 18 106 20 108
rect 26 106 28 108
rect 10 102 12 104
rect 18 102 20 104
rect 26 102 28 104
rect 10 98 12 100
rect 18 98 20 100
rect 26 98 28 100
rect 10 94 12 96
rect 18 94 20 96
rect 26 94 28 96
rect 14 73 16 75
rect 10 29 12 31
rect 18 29 20 31
rect 26 29 28 31
rect 10 25 12 27
rect 18 25 20 27
rect 26 25 28 27
rect 10 21 12 23
rect 18 21 20 23
rect 26 21 28 23
rect 10 17 12 19
rect 18 17 20 19
rect 26 17 28 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
rect 28 6 30 8
rect 32 6 34 8
<< poly >>
rect 14 91 16 128
rect 22 91 24 128
rect 14 89 24 91
rect 14 77 16 89
rect 12 71 18 77
rect 14 36 16 71
rect 14 34 24 36
rect 14 13 16 34
rect 22 13 24 34
<< ndiff >>
rect 6 130 36 136
rect 8 15 30 33
<< pdiff >>
rect 8 92 30 126
rect 6 4 36 10
<< nwell >>
rect 3 48 39 139
<< pwell >>
rect 3 1 39 46
<< end >>
