magic
tech concept
timestamp 1576254708844
<< metal1 >>
rect 0 133 28 138
rect 0 131 7 133
rect 9 131 12 133
rect 14 131 17 133
rect 19 131 28 133
rect 0 127 28 131
rect 8 123 12 127
rect 16 123 20 124
rect 8 121 9 123
rect 11 121 12 123
rect 16 121 17 123
rect 19 121 20 123
rect 8 119 12 121
rect 16 119 20 121
rect 8 117 9 119
rect 11 117 12 119
rect 16 117 17 119
rect 19 117 20 119
rect 8 115 12 117
rect 16 115 20 117
rect 8 113 9 115
rect 11 113 12 115
rect 16 113 17 115
rect 19 113 20 115
rect 8 111 12 113
rect 16 111 20 113
rect 8 109 9 111
rect 11 109 12 111
rect 16 109 17 111
rect 19 109 20 111
rect 8 107 12 109
rect 16 107 20 109
rect 8 105 9 107
rect 11 105 12 107
rect 16 105 17 107
rect 19 105 20 107
rect 8 103 12 105
rect 16 103 20 105
rect 8 101 9 103
rect 11 101 12 103
rect 16 101 17 103
rect 19 101 20 103
rect 8 99 12 101
rect 16 99 20 101
rect 8 97 9 99
rect 11 97 12 99
rect 16 97 17 99
rect 19 97 20 99
rect 8 95 12 97
rect 16 95 20 97
rect 8 93 9 95
rect 11 93 12 95
rect 16 93 17 95
rect 19 93 20 95
rect 8 92 12 93
rect 16 75 20 93
rect 8 66 12 75
rect 16 71 26 75
rect 16 30 20 71
rect 8 64 9 66
rect 11 64 12 66
rect 8 63 12 64
rect 8 30 12 31
rect 8 28 9 30
rect 11 28 12 30
rect 16 28 17 30
rect 19 28 20 30
rect 8 26 12 28
rect 16 26 20 28
rect 8 24 9 26
rect 11 24 12 26
rect 16 24 17 26
rect 19 24 20 26
rect 8 22 12 24
rect 16 22 20 24
rect 8 20 9 22
rect 11 20 12 22
rect 16 20 17 22
rect 19 20 20 22
rect 8 18 12 20
rect 16 18 20 20
rect 8 16 9 18
rect 11 16 12 18
rect 16 16 17 18
rect 19 16 20 18
rect 8 12 12 16
rect 16 15 20 16
rect 0 7 28 12
rect 0 5 7 7
rect 9 5 12 7
rect 14 5 17 7
rect 19 5 28 7
rect 0 1 28 5
<< contact >>
rect 7 131 9 133
rect 12 131 14 133
rect 17 131 19 133
rect 9 121 11 123
rect 17 121 19 123
rect 9 117 11 119
rect 17 117 19 119
rect 9 113 11 115
rect 17 113 19 115
rect 9 109 11 111
rect 17 109 19 111
rect 9 105 11 107
rect 17 105 19 107
rect 9 101 11 103
rect 17 101 19 103
rect 9 97 11 99
rect 17 97 19 99
rect 9 93 11 95
rect 17 93 19 95
rect 9 64 11 66
rect 9 28 11 30
rect 17 28 19 30
rect 9 24 11 26
rect 17 24 19 26
rect 9 20 11 22
rect 17 20 19 22
rect 9 16 11 18
rect 17 16 19 18
rect 7 5 9 7
rect 12 5 14 7
rect 17 5 19 7
<< poly >>
rect 13 68 15 127
rect 7 62 15 68
rect 13 12 15 62
<< ndiff >>
rect 5 129 23 135
rect 7 14 21 32
<< pdiff >>
rect 7 91 21 125
rect 5 3 23 9
<< nwell >>
rect 2 47 26 138
<< pwell >>
rect 2 0 26 45
<< end >>
