magic
tech concept
timestamp 1577734651598
<< sizer >>
rect 0 0 56 70
<< metal1 >>
rect 0 65 56 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 45 65
rect 47 63 49 65
rect 51 63 56 65
rect 0 58 56 63
rect 6 55 10 58
rect 35 55 39 58
rect 26 55 30 56
rect 43 55 47 56
rect 6 53 7 55
rect 9 53 10 55
rect 26 53 27 55
rect 29 53 30 55
rect 35 53 36 55
rect 38 53 39 55
rect 43 53 44 55
rect 46 53 47 55
rect 6 51 10 53
rect 26 51 30 53
rect 35 51 39 53
rect 43 51 47 53
rect 6 49 7 51
rect 9 49 10 51
rect 26 49 27 51
rect 29 49 30 51
rect 35 49 36 51
rect 38 49 39 51
rect 43 49 44 51
rect 46 49 53 51
rect 6 48 10 49
rect 26 48 30 49
rect 35 48 39 49
rect 43 48 53 49
rect 27 39 30 48
rect 50 41 53 48
rect 39 44 43 45
rect 39 42 40 44
rect 42 42 43 44
rect 39 41 43 42
rect 39 39 42 41
rect 50 37 54 41
rect 27 36 45 39
rect 50 19 53 37
rect 42 26 45 36
rect 1 33 12 34
rect 15 32 20 34
rect 22 32 28 34
rect 32 33 40 34
rect 1 31 9 33
rect 11 31 12 33
rect 32 31 33 33
rect 35 31 40 33
rect 15 30 17 32
rect 19 30 20 32
rect 22 30 25 32
rect 27 30 28 32
rect 1 30 5 31
rect 8 30 12 31
rect 32 30 40 31
rect 15 29 20 30
rect 24 29 28 30
rect 42 25 46 26
rect 42 24 43 25
rect 45 23 46 25
rect 15 23 43 24
rect 15 21 46 23
rect 15 19 18 21
rect 30 19 33 21
rect 6 18 10 19
rect 14 18 18 19
rect 22 18 26 19
rect 30 18 34 19
rect 38 18 42 19
rect 46 18 53 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 30 16 31 18
rect 33 16 34 18
rect 38 16 39 18
rect 41 16 42 18
rect 46 16 47 18
rect 49 16 53 18
rect 6 13 10 16
rect 14 15 18 16
rect 22 13 26 16
rect 30 15 34 16
rect 38 13 42 16
rect 46 15 53 16
rect 0 7 56 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 45 7
rect 47 5 49 7
rect 51 5 56 7
rect 0 2 56 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 45 63 47 65
rect 49 63 51 65
rect 7 53 9 55
rect 27 53 29 55
rect 36 53 38 55
rect 44 53 46 55
rect 7 49 9 51
rect 27 49 29 51
rect 36 49 38 51
rect 44 49 46 51
rect 40 42 42 44
rect 9 31 11 33
rect 33 31 35 33
rect 17 30 19 32
rect 25 30 27 32
rect 43 23 45 25
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 31 16 33 18
rect 39 16 41 18
rect 47 16 49 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
rect 45 5 47 7
rect 49 5 51 7
<< poly >>
rect 11 35 13 59
rect 15 34 17 59
rect 19 38 21 59
rect 23 42 25 59
rect 40 46 42 59
rect 38 40 44 46
rect 23 40 33 42
rect 31 35 33 40
rect 19 36 25 38
rect 23 34 25 36
rect 7 29 13 35
rect 31 29 37 35
rect 15 28 21 34
rect 23 28 29 34
rect 11 12 13 29
rect 35 12 37 29
rect 19 12 21 28
rect 27 12 29 28
rect 41 21 47 27
rect 43 12 45 21
<< ndiff >>
rect 3 61 53 67
rect 5 14 51 20
<< pdiff >>
rect 5 47 31 57
rect 34 47 48 57
rect 3 3 53 9
<< nwell >>
rect 0 31 56 70
<< pwell >>
rect 0 0 56 31
<< end >>
