magic
tech scmos
timestamp 1573846977975
<< nwell >>
rect 9 196 45 212
<< pwell >>
rect 10 171 40 185
<< polysilicon >>
rect 21 203 24 204
rect 29 203 32 204
rect 21 196 24 198
rect 29 190 32 198
rect 10 196 15 197
rect 10 193 11 196
rect 14 193 24 196
rect 10 192 15 193
rect 21 183 24 193
rect 28 189 33 190
rect 28 186 29 189
rect 32 186 33 189
rect 28 185 33 186
rect 29 183 32 185
rect 21 177 24 178
rect 29 177 32 178
<< ndiffusion >>
rect 15 182 21 183
rect 24 178 29 183
rect 32 182 38 183
rect 15 179 16 182
rect 19 179 21 182
rect 32 179 34 182
rect 37 179 38 182
rect 15 178 21 179
rect 32 178 38 179
<< pdiffusion >>
rect 15 209 20 210
rect 33 209 38 210
rect 15 206 16 209
rect 19 206 20 209
rect 33 206 34 209
rect 37 206 38 209
rect 15 203 20 206
rect 33 203 38 206
rect 15 198 21 203
rect 24 202 29 203
rect 32 198 38 203
rect 24 199 25 202
rect 28 199 29 202
rect 24 198 29 199
<< ntransistor >>
rect 21 178 24 183
rect 29 178 32 183
<< ptransistor >>
rect 21 198 24 203
rect 29 198 32 203
<< polycontact >>
rect 11 193 14 196
rect 29 186 32 189
<< ndcontact >>
rect 16 179 19 182
rect 34 179 37 182
<< pdcontact >>
rect 16 206 19 209
rect 34 206 37 209
rect 25 199 28 202
<< nsubstratencontact >>
rect 11 206 14 209
rect 22 206 25 209
rect 28 206 31 209
rect 40 206 43 209
<< psubstratepcontact >>
rect 11 172 14 175
rect 16 172 19 175
rect 21 172 24 175
rect 26 172 29 175
rect 31 172 34 175
rect 36 172 39 175
<< metal1 >>
rect 0 205 47 210
rect 24 197 29 203
rect 0 192 15 197
rect 24 192 40 197
rect 35 187 47 192
rect 0 185 33 190
rect 35 183 40 187
rect 15 176 20 183
rect 33 178 40 183
rect 0 171 47 176
<< labels >>
rlabel metal1 0 205 47 210 1 vdd
rlabel metal1 0 171 47 176 1 gnd
rlabel metal1 0 192 15 197 1 inX
rlabel metal1 0 185 33 190 1 inY
rlabel metal1 35 187 47 192 1 out
<< end >>
