magic
tech concept
timestamp 1576599475403
<< sizer >>
rect 0 0 42 140
<< metal1 >>
rect 0 134 42 139
rect 0 132 8 134
rect 10 132 12 134
rect 14 132 16 134
rect 18 132 20 134
rect 22 132 24 134
rect 26 132 28 134
rect 30 132 32 134
rect 34 132 42 134
rect 0 128 42 132
rect 17 124 21 128
rect 31 109 34 128
rect 9 124 13 125
rect 25 124 29 125
rect 9 122 10 124
rect 12 122 13 124
rect 17 122 18 124
rect 20 122 21 124
rect 25 122 26 124
rect 28 122 29 124
rect 9 120 13 122
rect 17 120 21 122
rect 25 120 29 122
rect 9 118 10 120
rect 12 118 13 120
rect 17 118 18 120
rect 20 118 21 120
rect 25 118 26 120
rect 28 118 29 120
rect 9 115 13 118
rect 17 117 21 118
rect 25 115 29 118
rect 2 116 6 117
rect 2 114 3 116
rect 5 114 6 116
rect 9 111 29 115
rect 2 113 6 114
rect 2 90 5 113
rect 14 49 17 111
rect 8 108 12 109
rect 22 106 34 109
rect 8 106 9 108
rect 11 106 12 108
rect 8 105 12 106
rect 22 62 25 106
rect 8 76 11 105
rect 1 86 5 90
rect 2 27 5 86
rect 8 72 12 76
rect 8 35 11 72
rect 21 61 25 62
rect 29 61 33 62
rect 21 59 22 61
rect 24 59 25 61
rect 29 59 30 61
rect 32 59 33 61
rect 21 57 25 59
rect 29 57 33 59
rect 21 55 22 57
rect 24 55 25 57
rect 29 55 30 57
rect 32 55 33 57
rect 21 54 25 55
rect 29 54 33 55
rect 30 40 33 54
rect 14 48 23 49
rect 14 46 20 48
rect 22 46 23 48
rect 19 45 23 46
rect 20 20 23 45
rect 36 40 40 41
rect 29 39 40 40
rect 29 37 30 39
rect 32 37 40 39
rect 29 36 33 37
rect 8 34 12 35
rect 8 32 9 34
rect 11 32 12 34
rect 8 31 12 32
rect 29 31 33 32
rect 29 29 30 31
rect 32 29 33 31
rect 29 28 33 29
rect 30 13 33 28
rect 2 26 7 27
rect 2 24 4 26
rect 6 24 7 26
rect 2 23 7 24
rect 9 19 13 20
rect 20 19 25 20
rect 9 17 10 19
rect 12 17 13 19
rect 20 17 22 19
rect 24 17 25 19
rect 9 13 13 17
rect 20 16 25 17
rect 0 8 42 13
rect 0 6 8 8
rect 10 6 12 8
rect 14 6 16 8
rect 18 6 20 8
rect 22 6 24 8
rect 26 6 28 8
rect 30 6 32 8
rect 34 6 42 8
rect 0 2 42 6
<< contact >>
rect 8 132 10 134
rect 12 132 14 134
rect 16 132 18 134
rect 20 132 22 134
rect 24 132 26 134
rect 28 132 30 134
rect 32 132 34 134
rect 10 122 12 124
rect 18 122 20 124
rect 26 122 28 124
rect 10 118 12 120
rect 18 118 20 120
rect 26 118 28 120
rect 3 114 5 116
rect 9 106 11 108
rect 22 59 24 61
rect 30 59 32 61
rect 22 55 24 57
rect 30 55 32 57
rect 20 46 22 48
rect 30 37 32 39
rect 9 32 11 34
rect 30 29 32 31
rect 4 24 6 26
rect 10 17 12 19
rect 22 17 24 19
rect 8 6 10 8
rect 12 6 14 8
rect 16 6 18 8
rect 20 6 22 8
rect 24 6 26 8
rect 28 6 30 8
rect 32 6 34 8
<< poly >>
rect 14 115 16 128
rect 22 110 24 128
rect 1 115 7 118
rect 1 113 16 115
rect 1 112 7 113
rect 7 108 24 110
rect 7 104 13 108
rect 26 50 28 65
rect 18 48 28 50
rect 18 44 24 48
rect 21 35 23 44
rect 7 30 13 36
rect 21 33 36 35
rect 10 28 12 30
rect 2 24 8 28
rect 10 26 20 28
rect 18 13 20 26
rect 2 22 16 24
rect 14 13 16 22
<< ndiff >>
rect 6 130 36 136
rect 28 27 34 41
rect 8 15 26 21
<< pdiff >>
rect 8 116 30 126
rect 20 53 34 63
rect 6 4 36 10
<< nwell >>
rect 3 48 39 139
<< pwell >>
rect 3 1 39 46
<< end >>
