magic
tech concept
timestamp 1577797116938
<< sizer >>
rect 0 0 42 70
<< metal1 >>
rect 0 65 42 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 42 65
rect 0 58 42 63
rect 6 55 14 58
rect 28 55 36 58
rect 6 53 7 55
rect 9 53 11 55
rect 13 53 14 55
rect 28 53 29 55
rect 31 53 33 55
rect 35 53 36 55
rect 6 52 14 53
rect 28 52 36 53
rect 6 47 14 48
rect 6 45 7 47
rect 9 45 11 47
rect 13 45 14 47
rect 6 44 14 45
rect 8 41 11 44
rect 28 43 36 44
rect 28 41 29 43
rect 31 41 33 43
rect 35 41 39 43
rect 2 40 6 41
rect 8 40 14 41
rect 28 40 39 41
rect 2 38 3 40
rect 5 38 6 40
rect 8 38 11 40
rect 13 38 14 40
rect 36 34 39 40
rect 2 37 6 38
rect 8 37 14 38
rect 8 26 11 37
rect 22 33 26 34
rect 36 30 40 34
rect 22 31 23 33
rect 25 31 26 33
rect 22 30 26 31
rect 36 19 39 30
rect 7 25 11 26
rect 7 23 8 25
rect 10 23 11 25
rect 7 22 11 23
rect 17 18 21 19
rect 29 18 39 19
rect 7 17 11 18
rect 17 16 18 18
rect 20 16 21 18
rect 29 16 30 18
rect 32 16 39 18
rect 7 15 8 17
rect 10 15 11 17
rect 17 13 21 16
rect 29 15 33 16
rect 7 13 11 15
rect 0 7 42 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 42 7
rect 0 2 42 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 7 53 9 55
rect 11 53 13 55
rect 29 53 31 55
rect 33 53 35 55
rect 7 45 9 47
rect 11 45 13 47
rect 29 41 31 43
rect 33 41 35 43
rect 3 38 5 40
rect 11 38 13 40
rect 23 31 25 33
rect 8 23 10 25
rect 18 16 20 18
rect 30 16 32 18
rect 8 15 10 17
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
<< poly >>
rect 2 49 17 51
rect 19 49 39 51
rect 2 42 4 49
rect 19 47 21 49
rect 16 45 21 47
rect 23 45 39 47
rect 16 42 18 45
rect 23 35 25 45
rect 1 36 7 42
rect 9 40 18 42
rect 9 36 15 40
rect 2 21 4 36
rect 21 32 27 35
rect 21 29 28 32
rect 26 12 28 29
rect 13 21 24 23
rect 2 19 15 21
rect 22 12 24 21
<< ndiff >>
rect 3 61 39 67
rect 6 13 12 27
rect 16 14 34 20
<< pdiff >>
rect 5 43 15 57
rect 27 39 37 57
rect 3 3 39 9
<< nwell >>
rect 0 32 42 70
rect 17 31 42 32
<< pwell >>
rect 0 31 17 32
rect 0 0 42 31
<< end >>
