magic
tech concept
timestamp 1577134497824
<< sizer >>
rect 0 0 35 70
<< metal1 >>
rect 0 65 35 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 35 65
rect 0 58 35 63
rect 14 55 18 58
rect 6 55 10 56
rect 22 55 26 56
rect 6 53 7 55
rect 9 53 10 55
rect 14 53 15 55
rect 17 53 18 55
rect 22 53 23 55
rect 25 53 26 55
rect 6 51 10 53
rect 14 51 18 53
rect 22 51 26 53
rect 6 49 7 51
rect 9 49 12 51
rect 14 49 15 51
rect 17 49 18 51
rect 22 49 23 51
rect 25 49 26 51
rect 6 48 12 49
rect 14 48 18 49
rect 22 48 26 49
rect 9 33 12 48
rect 23 34 26 48
rect 1 33 6 34
rect 23 31 33 34
rect 1 31 3 33
rect 5 31 6 33
rect 9 32 20 33
rect 9 30 17 32
rect 19 30 20 32
rect 1 30 6 31
rect 23 19 26 31
rect 29 30 33 31
rect 9 29 20 30
rect 9 19 12 29
rect 6 18 12 19
rect 14 18 18 19
rect 22 18 26 19
rect 6 16 7 18
rect 9 16 12 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 6 15 12 16
rect 14 13 18 16
rect 22 15 26 16
rect 0 7 35 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 35 7
rect 0 2 35 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 7 53 9 55
rect 15 53 17 55
rect 23 53 25 55
rect 7 49 9 51
rect 15 49 17 51
rect 23 49 25 51
rect 3 31 5 33
rect 17 30 19 32
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
<< poly >>
rect 11 46 13 59
rect 19 34 21 59
rect 5 44 13 46
rect 5 35 7 44
rect 1 29 7 35
rect 15 28 21 34
rect 5 23 7 29
rect 19 12 21 28
rect 5 21 13 23
rect 11 12 13 21
<< ndiff >>
rect 3 61 29 67
rect 5 14 27 20
<< pdiff >>
rect 5 47 27 57
rect 3 3 25 9
<< nwell >>
rect 0 31 35 70
<< pwell >>
rect 0 0 35 31
<< end >>
