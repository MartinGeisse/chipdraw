magic
tech concept
timestamp 1577188023699
<< sizer >>
rect 0 0 42 70
<< metal1 >>
rect 0 65 42 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 42 65
rect 0 58 42 63
rect 6 55 10 58
rect 22 55 26 56
rect 6 53 7 55
rect 9 53 10 55
rect 22 53 23 55
rect 25 53 26 55
rect 6 51 10 53
rect 22 51 26 53
rect 6 49 7 51
rect 9 49 10 51
rect 15 49 23 51
rect 25 49 26 51
rect 6 48 10 49
rect 15 48 26 49
rect 15 34 18 48
rect 1 33 12 34
rect 15 30 19 34
rect 22 33 26 34
rect 29 33 34 34
rect 1 31 9 33
rect 11 31 12 33
rect 22 31 23 33
rect 25 31 26 33
rect 29 31 31 33
rect 33 31 34 33
rect 1 30 5 31
rect 8 30 12 31
rect 22 30 26 31
rect 29 30 34 31
rect 15 24 18 30
rect 15 21 33 24
rect 15 19 18 21
rect 30 19 33 21
rect 6 18 10 19
rect 14 18 18 19
rect 22 18 26 19
rect 30 18 34 19
rect 6 16 7 18
rect 9 16 10 18
rect 14 16 15 18
rect 17 16 18 18
rect 22 16 23 18
rect 25 16 26 18
rect 30 16 31 18
rect 33 16 34 18
rect 6 13 10 16
rect 14 15 18 16
rect 22 13 26 16
rect 30 15 34 16
rect 0 7 42 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 34 7
rect 36 5 42 7
rect 0 2 42 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 7 53 9 55
rect 23 53 25 55
rect 7 49 9 51
rect 23 49 25 51
rect 9 31 11 33
rect 23 31 25 33
rect 31 31 33 33
rect 7 16 9 18
rect 15 16 17 18
rect 23 16 25 18
rect 31 16 33 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 34 5 36 7
<< poly >>
rect 11 35 13 59
rect 15 35 17 59
rect 19 42 21 59
rect 19 40 31 42
rect 29 35 31 40
rect 7 29 13 35
rect 15 33 27 35
rect 29 29 35 35
rect 19 29 27 33
rect 11 12 13 29
rect 19 12 21 29
rect 29 25 31 29
rect 27 23 31 25
rect 27 12 29 23
<< ndiff >>
rect 3 61 37 67
rect 5 14 35 20
<< pdiff >>
rect 5 47 27 57
rect 3 3 38 9
<< nwell >>
rect 0 31 42 70
<< pwell >>
rect 0 0 42 31
<< end >>
