magic
tech LibreSilicon-test000-concept-mg-70-7
timestamp 1577186511752
<< sizer >>
rect 0 0 49 70
<< metal1 >>
rect 0 65 49 69
rect 0 63 5 65
rect 7 63 9 65
rect 11 63 13 65
rect 15 63 17 65
rect 19 63 21 65
rect 23 63 25 65
rect 27 63 29 65
rect 31 63 33 65
rect 35 63 37 65
rect 39 63 41 65
rect 43 63 49 65
rect 0 58 49 63
rect 14 50 18 58
rect 22 53 42 56
rect 22 50 26 53
rect 38 50 42 53
rect 6 50 10 51
rect 30 50 34 51
rect 6 48 7 50
rect 9 48 10 50
rect 14 48 15 50
rect 17 48 18 50
rect 22 48 23 50
rect 25 48 26 50
rect 30 48 31 50
rect 33 48 34 50
rect 38 48 39 50
rect 41 48 42 50
rect 6 46 10 48
rect 14 46 18 48
rect 22 46 26 48
rect 30 46 34 48
rect 38 46 42 48
rect 6 44 7 46
rect 9 44 10 46
rect 14 44 15 46
rect 17 44 18 46
rect 22 44 23 46
rect 25 44 26 46
rect 30 44 31 46
rect 33 44 34 46
rect 38 44 39 46
rect 41 44 42 46
rect 6 41 10 44
rect 14 43 18 44
rect 22 41 26 44
rect 30 43 34 44
rect 38 43 42 44
rect 31 41 34 43
rect 6 38 26 41
rect 31 38 46 41
rect 43 34 46 38
rect 8 33 12 34
rect 15 33 20 34
rect 29 33 33 34
rect 36 33 41 34
rect 43 30 47 34
rect 8 31 9 33
rect 11 31 12 33
rect 15 31 17 33
rect 19 31 20 33
rect 29 31 30 33
rect 32 31 33 33
rect 36 31 38 33
rect 40 31 41 33
rect 8 30 12 31
rect 15 30 20 31
rect 29 30 33 31
rect 36 30 41 31
rect 43 24 46 30
rect 19 21 46 24
rect 19 19 22 21
rect 6 18 10 19
rect 18 18 22 19
rect 30 18 34 19
rect 6 16 7 18
rect 9 16 10 18
rect 18 16 19 18
rect 21 16 22 18
rect 30 16 31 18
rect 33 16 34 18
rect 6 13 10 16
rect 18 15 22 16
rect 30 13 34 16
rect 0 7 49 13
rect 0 5 5 7
rect 7 5 9 7
rect 11 5 13 7
rect 15 5 17 7
rect 19 5 21 7
rect 23 5 25 7
rect 27 5 29 7
rect 31 5 33 7
rect 35 5 37 7
rect 39 5 41 7
rect 43 5 49 7
rect 0 2 49 5
<< contact >>
rect 5 63 7 65
rect 9 63 11 65
rect 13 63 15 65
rect 17 63 19 65
rect 21 63 23 65
rect 25 63 27 65
rect 29 63 31 65
rect 33 63 35 65
rect 37 63 39 65
rect 41 63 43 65
rect 7 48 9 50
rect 15 48 17 50
rect 23 48 25 50
rect 31 48 33 50
rect 39 48 41 50
rect 7 44 9 46
rect 15 44 17 46
rect 23 44 25 46
rect 31 44 33 46
rect 39 44 41 46
rect 9 31 11 33
rect 17 31 19 33
rect 30 31 32 33
rect 38 31 40 33
rect 7 16 9 18
rect 19 16 21 18
rect 31 16 33 18
rect 5 5 7 7
rect 9 5 11 7
rect 13 5 15 7
rect 17 5 19 7
rect 21 5 23 7
rect 25 5 27 7
rect 29 5 31 7
rect 33 5 35 7
rect 37 5 39 7
rect 41 5 43 7
<< poly >>
rect 11 35 13 54
rect 19 35 21 54
rect 27 41 29 54
rect 35 41 37 54
rect 27 39 30 41
rect 35 39 38 41
rect 28 35 30 39
rect 36 35 38 39
rect 7 29 13 35
rect 15 29 21 35
rect 28 29 34 35
rect 36 29 42 35
rect 11 12 13 29
rect 15 12 17 29
rect 28 27 30 29
rect 36 23 38 29
rect 23 25 30 27
rect 23 12 25 25
rect 27 21 38 23
rect 27 12 29 21
<< ndiff >>
rect 3 61 45 67
rect 5 14 35 20
<< pdiff >>
rect 5 42 43 52
rect 3 3 45 9
<< nwell >>
rect 0 31 49 70
<< pwell >>
rect 0 0 49 31
<< end >>
